magic
tech sky130A
magscale 1 2
timestamp 1666517498
<< error_s >>
rect 1352 -1136 1474 -1133
rect 1380 -1164 1446 -1161
rect 1387 -1175 1439 -1168
<< locali >>
rect -81 244 -16 259
rect -81 208 -66 244
rect -30 208 -16 244
rect 274 246 330 261
rect -81 193 -16 208
rect 274 210 284 246
rect 320 210 330 246
rect 1843 256 1909 265
rect 1843 220 1858 256
rect 1894 220 1909 256
rect 1843 211 1909 220
rect 2013 256 2079 265
rect 2013 220 2028 256
rect 2064 220 2079 256
rect 2013 211 2079 220
rect 274 195 330 210
rect 1937 119 1985 125
rect 1937 85 1944 119
rect 1978 85 1985 119
rect 1937 78 1985 85
rect 1380 -129 1446 -114
rect 1380 -165 1395 -129
rect 1431 -165 1446 -129
rect 1421 -180 1446 -165
rect 274 -210 330 -195
rect 274 -246 284 -210
rect 320 -246 330 -210
rect 274 -261 330 -246
rect 274 -842 330 -827
rect 274 -878 284 -842
rect 320 -878 330 -842
rect 274 -893 330 -878
rect 1422 -923 1446 -908
rect 1380 -959 1395 -923
rect 1431 -959 1446 -923
rect 1380 -974 1446 -959
rect 1385 -1183 1441 -1168
rect 1385 -1219 1395 -1183
rect 1431 -1219 1441 -1183
rect 1385 -1234 1441 -1219
rect 1944 -1206 1998 -1191
rect 1944 -1242 1952 -1206
rect 1988 -1242 1998 -1206
rect 1944 -1257 1998 -1242
rect 1944 -1258 1994 -1257
rect 16 -1299 82 -1284
rect 16 -1335 31 -1299
rect 67 -1335 82 -1299
rect 16 -1350 82 -1335
rect 275 -1301 329 -1286
rect 275 -1337 283 -1301
rect 319 -1337 329 -1301
rect 275 -1352 329 -1337
rect 2012 -1309 2078 -1299
rect 2012 -1345 2027 -1309
rect 2063 -1345 2078 -1309
rect 275 -1353 325 -1352
rect 2012 -1353 2078 -1345
rect 1669 -1837 1735 -1822
rect 1669 -1873 1684 -1837
rect 1720 -1873 1735 -1837
rect 1711 -1888 1735 -1873
rect 18 -1914 88 -1913
rect 16 -1929 88 -1914
rect 16 -1965 31 -1929
rect 67 -1965 88 -1929
rect 16 -1980 88 -1965
rect 274 -1930 330 -1920
rect 274 -1966 284 -1930
rect 320 -1966 330 -1930
rect 274 -1976 330 -1966
rect 1385 -2045 1441 -2030
rect 1385 -2081 1395 -2045
rect 1431 -2081 1441 -2045
rect 1385 -2096 1441 -2081
<< viali >>
rect -66 208 -30 244
rect 29 212 69 252
rect 284 210 320 246
rect 1858 220 1894 256
rect 2028 220 2064 256
rect 1395 129 1431 165
rect 1944 85 1978 119
rect 1395 -165 1431 -129
rect 29 -252 69 -212
rect 284 -246 320 -210
rect 29 -876 69 -836
rect 284 -878 320 -842
rect 1395 -959 1431 -923
rect 1395 -1219 1431 -1183
rect 1952 -1242 1988 -1206
rect 31 -1335 67 -1299
rect 283 -1337 319 -1301
rect 1860 -1346 1900 -1306
rect 2027 -1345 2063 -1309
rect 1684 -1873 1720 -1837
rect 31 -1965 67 -1929
rect 284 -1966 320 -1930
rect 1395 -2081 1431 -2045
<< metal1 >>
rect 1748 496 1824 592
rect -81 252 -16 259
rect 22 252 78 265
rect 1843 264 1909 271
rect -81 200 -74 252
rect -22 212 29 252
rect 69 212 78 252
rect -22 200 78 212
rect -81 199 78 200
rect 269 254 335 261
rect 269 202 276 254
rect 328 248 335 254
rect 328 208 1528 248
rect 328 202 335 208
rect -81 193 -16 199
rect 269 195 335 202
rect -68 -199 -28 193
rect 1380 173 1446 180
rect 1380 121 1387 173
rect 1439 121 1446 173
rect 1380 114 1446 121
rect 1488 122 1528 208
rect 1843 212 1850 264
rect 1902 212 1909 264
rect 1843 205 1909 212
rect 2013 264 2079 271
rect 2013 212 2020 264
rect 2072 212 2079 264
rect 2013 205 2079 212
rect 1932 122 1990 131
rect 1488 119 1990 122
rect 1488 85 1944 119
rect 1978 85 1990 119
rect 1488 82 1990 85
rect 1932 76 1990 82
rect 1748 -48 1824 48
rect 1380 -121 1446 -114
rect 1380 -173 1387 -121
rect 1439 -127 1446 -121
rect 1844 -127 1850 -121
rect 1439 -167 1850 -127
rect 1439 -173 1446 -167
rect 1844 -173 1850 -167
rect 1902 -173 1908 -121
rect 1380 -180 1446 -173
rect -68 -212 78 -199
rect -68 -252 29 -212
rect 69 -252 78 -212
rect -68 -265 78 -252
rect 269 -202 335 -195
rect 269 -254 276 -202
rect 328 -254 335 -202
rect 269 -261 335 -254
rect -68 -823 -28 -265
rect -68 -836 78 -823
rect -68 -876 29 -836
rect 69 -876 78 -836
rect 22 -889 78 -876
rect 269 -834 335 -827
rect 269 -886 276 -834
rect 328 -886 335 -834
rect 269 -893 335 -886
rect 1380 -915 1446 -908
rect 1380 -967 1387 -915
rect 1439 -921 1446 -915
rect 2013 -921 2019 -915
rect 1439 -961 2019 -921
rect 1439 -967 1446 -961
rect 2013 -967 2019 -961
rect 2071 -967 2077 -915
rect 1380 -974 1446 -967
rect 1748 -1136 1824 -1040
rect 1380 -1174 1446 -1161
rect 1380 -1175 1897 -1174
rect 1380 -1220 1387 -1175
rect 1439 -1214 1897 -1175
rect 1439 -1220 1446 -1214
rect 1380 -1227 1446 -1220
rect 16 -1297 82 -1284
rect 146 -1297 152 -1291
rect 16 -1299 152 -1297
rect 16 -1335 31 -1299
rect 67 -1335 152 -1299
rect 16 -1337 152 -1335
rect 16 -1350 82 -1337
rect 146 -1343 152 -1337
rect 204 -1343 210 -1291
rect 275 -1299 329 -1286
rect 1857 -1287 1897 -1214
rect 1937 -1198 2003 -1191
rect 1937 -1250 1944 -1198
rect 1996 -1250 2003 -1198
rect 1937 -1257 2003 -1250
rect 1756 -1299 1762 -1293
rect 275 -1301 1762 -1299
rect 275 -1337 283 -1301
rect 319 -1337 1762 -1301
rect 275 -1339 1762 -1337
rect 275 -1352 329 -1339
rect 1756 -1345 1762 -1339
rect 1814 -1345 1820 -1293
rect 1848 -1306 1912 -1287
rect 1848 -1346 1860 -1306
rect 1900 -1346 1912 -1306
rect 1848 -1353 1912 -1346
rect 2012 -1301 2078 -1294
rect 2012 -1353 2019 -1301
rect 2071 -1353 2078 -1301
rect 2012 -1360 2078 -1353
rect 1748 -1680 1824 -1584
rect 1669 -1835 1735 -1822
rect 1669 -1837 2138 -1835
rect 1669 -1873 1684 -1837
rect 1720 -1873 2138 -1837
rect 1669 -1875 2138 -1873
rect 1669 -1888 1735 -1875
rect 16 -1927 82 -1914
rect 146 -1927 152 -1921
rect 16 -1929 152 -1927
rect 16 -1965 31 -1929
rect 67 -1965 152 -1929
rect 16 -1967 152 -1965
rect 16 -1980 82 -1967
rect 146 -1973 152 -1967
rect 204 -1973 210 -1921
rect 269 -1922 335 -1915
rect 269 -1974 276 -1922
rect 328 -1974 335 -1922
rect 269 -1981 335 -1974
rect 1380 -2037 1446 -2030
rect 1380 -2089 1387 -2037
rect 1439 -2043 1446 -2037
rect 2013 -2043 2019 -2037
rect 1439 -2083 2019 -2043
rect 1439 -2089 1446 -2083
rect 2013 -2089 2019 -2083
rect 2071 -2089 2077 -2037
rect 1380 -2096 1446 -2089
<< via1 >>
rect 20 518 72 570
rect -74 244 -22 252
rect -74 208 -66 244
rect -66 208 -30 244
rect -30 208 -22 244
rect -74 200 -22 208
rect 276 246 328 254
rect 276 210 284 246
rect 284 210 320 246
rect 320 210 328 246
rect 276 202 328 210
rect 1387 165 1439 173
rect 1387 129 1395 165
rect 1395 129 1431 165
rect 1431 129 1439 165
rect 1387 121 1439 129
rect 1850 256 1902 264
rect 1850 220 1858 256
rect 1858 220 1894 256
rect 1894 220 1902 256
rect 1850 212 1902 220
rect 2020 256 2072 264
rect 2020 220 2028 256
rect 2028 220 2064 256
rect 2064 220 2072 256
rect 2020 212 2072 220
rect 1676 -26 1728 26
rect 1387 -129 1439 -121
rect 1387 -165 1395 -129
rect 1395 -165 1431 -129
rect 1431 -165 1439 -129
rect 1387 -173 1439 -165
rect 1850 -173 1902 -121
rect 276 -210 328 -202
rect 276 -246 284 -210
rect 284 -246 320 -210
rect 320 -246 328 -210
rect 276 -254 328 -246
rect 20 -570 72 -518
rect 276 -842 328 -834
rect 276 -878 284 -842
rect 284 -878 320 -842
rect 320 -878 328 -842
rect 276 -886 328 -878
rect 1387 -923 1439 -915
rect 1387 -959 1395 -923
rect 1395 -959 1431 -923
rect 1431 -959 1439 -923
rect 1387 -967 1439 -959
rect 2019 -967 2071 -915
rect 1676 -1114 1728 -1062
rect 1387 -1183 1439 -1175
rect 1387 -1219 1395 -1183
rect 1395 -1219 1431 -1183
rect 1431 -1219 1439 -1183
rect 1387 -1220 1439 -1219
rect 152 -1343 204 -1291
rect 1944 -1206 1996 -1198
rect 1944 -1242 1952 -1206
rect 1952 -1242 1988 -1206
rect 1988 -1242 1996 -1206
rect 1944 -1250 1996 -1242
rect 1762 -1345 1814 -1293
rect 2019 -1309 2071 -1301
rect 2019 -1345 2027 -1309
rect 2027 -1345 2063 -1309
rect 2063 -1345 2071 -1309
rect 2019 -1353 2071 -1345
rect 20 -1658 72 -1606
rect 152 -1973 204 -1921
rect 276 -1930 328 -1922
rect 276 -1966 284 -1930
rect 284 -1966 320 -1930
rect 320 -1966 328 -1930
rect 276 -1974 328 -1966
rect 1387 -2045 1439 -2037
rect 1387 -2081 1395 -2045
rect 1395 -2081 1431 -2045
rect 1431 -2081 1439 -2045
rect 1387 -2089 1439 -2081
rect 2019 -2089 2071 -2037
rect 1676 -2202 1728 -2150
<< metal2 >>
rect 14 570 78 697
rect 14 518 20 570
rect 72 518 78 570
rect -81 252 -16 259
rect -81 200 -74 252
rect -22 200 -16 252
rect -81 193 -16 200
rect 14 -518 78 518
rect 269 254 335 261
rect 269 202 276 254
rect 328 202 335 254
rect 269 195 335 202
rect 1380 173 1446 180
rect 1380 167 1387 173
rect 282 127 1387 167
rect 282 -195 322 127
rect 1380 121 1387 127
rect 1439 121 1446 173
rect 1380 114 1446 121
rect 1670 26 1734 697
rect 1843 264 1909 271
rect 1843 212 1850 264
rect 1902 212 1909 264
rect 1843 205 1909 212
rect 2013 264 2079 271
rect 2013 212 2020 264
rect 2072 212 2079 264
rect 2013 205 2079 212
rect 1670 -26 1676 26
rect 1728 -26 1734 26
rect 1380 -121 1446 -114
rect 1380 -173 1387 -121
rect 1439 -173 1446 -121
rect 1380 -180 1446 -173
rect 269 -202 335 -195
rect 269 -208 276 -202
rect 14 -570 20 -518
rect 72 -570 78 -518
rect 14 -1606 78 -570
rect 158 -248 276 -208
rect 158 -1285 198 -248
rect 269 -254 276 -248
rect 328 -254 335 -202
rect 269 -261 335 -254
rect 269 -834 335 -827
rect 269 -886 276 -834
rect 328 -840 335 -834
rect 1393 -840 1433 -180
rect 328 -880 1433 -840
rect 328 -886 335 -880
rect 269 -893 335 -886
rect 1380 -915 1446 -908
rect 1380 -967 1387 -915
rect 1439 -967 1446 -915
rect 1380 -974 1446 -967
rect 1670 -1062 1734 -26
rect 1856 -115 1896 205
rect 1850 -121 1902 -115
rect 1850 -179 1902 -173
rect 2025 -909 2065 205
rect 2019 -915 2071 -909
rect 2019 -973 2071 -967
rect 1670 -1114 1676 -1062
rect 1728 -1114 1734 -1062
rect 1380 -1175 1446 -1168
rect 1380 -1181 1387 -1175
rect 282 -1220 1387 -1181
rect 1439 -1220 1446 -1175
rect 282 -1221 1446 -1220
rect 152 -1291 204 -1285
rect 152 -1349 204 -1343
rect 14 -1658 20 -1606
rect 72 -1658 78 -1606
rect 14 -1665 78 -1658
rect 158 -1915 198 -1349
rect 282 -1915 322 -1221
rect 1380 -1234 1446 -1221
rect 152 -1921 204 -1915
rect 152 -1979 204 -1973
rect 269 -1922 335 -1915
rect 269 -1974 276 -1922
rect 328 -1974 335 -1922
rect 158 -1994 198 -1979
rect 269 -1981 335 -1974
rect 1380 -2037 1446 -2030
rect 1380 -2089 1387 -2037
rect 1439 -2089 1446 -2037
rect 1380 -2096 1446 -2089
rect 1670 -2150 1734 -1114
rect 1937 -1198 2003 -1191
rect 1937 -1204 1944 -1198
rect 1768 -1244 1944 -1204
rect 1768 -1287 1808 -1244
rect 1937 -1250 1944 -1244
rect 1996 -1250 2003 -1198
rect 1937 -1257 2003 -1250
rect 1762 -1293 1814 -1287
rect 1762 -1351 1814 -1345
rect 2012 -1301 2078 -1294
rect 2012 -1353 2019 -1301
rect 2071 -1353 2078 -1301
rect 2012 -1360 2078 -1353
rect 2025 -2031 2065 -1360
rect 2019 -2037 2071 -2031
rect 2019 -2095 2071 -2089
rect 1670 -2202 1676 -2150
rect 1728 -2202 1734 -2150
rect 1670 -2224 1734 -2202
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 0 0 1 0
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_1
timestamp 1644511149
transform 1 0 0 0 -1 0
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_2
timestamp 1644511149
transform 1 0 0 0 1 -1088
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_3
timestamp 1644511149
transform 1 0 0 0 -1 -1088
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_4
timestamp 1644511149
transform 1 0 0 0 1 -2176
box -38 -48 1786 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1824 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_1
timestamp 1644511149
transform 1 0 1824 0 -1 -1088
box -38 -48 314 592
<< labels >>
rlabel metal1 -68 -265 -2 -199 0 clk_in
rlabel metal2 14 633 78 697 0 vdd
rlabel metal2 1670 633 1734 697 5 vss
rlabel metal1 2098 -1875 2138 -1835 7 clk_out
<< end >>
