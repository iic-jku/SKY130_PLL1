magic
tech sky130A
magscale 1 2
timestamp 1652802024
<< nwell >>
rect -359 -289 359 289
<< pmos >>
rect -159 -70 -129 70
rect -63 -70 -33 70
rect 33 -70 63 70
rect 129 -70 159 70
<< pdiff >>
rect -221 58 -159 70
rect -221 -58 -209 58
rect -175 -58 -159 58
rect -221 -70 -159 -58
rect -129 58 -63 70
rect -129 -58 -113 58
rect -79 -58 -63 58
rect -129 -70 -63 -58
rect -33 58 33 70
rect -33 -58 -17 58
rect 17 -58 33 58
rect -33 -70 33 -58
rect 63 58 129 70
rect 63 -58 79 58
rect 113 -58 129 58
rect 63 -70 129 -58
rect 159 58 225 70
rect 159 -58 175 58
rect 209 -58 225 58
rect 159 -70 225 -58
<< pdiffc >>
rect -209 -58 -175 58
rect -113 -58 -79 58
rect -17 -58 17 58
rect 79 -58 113 58
rect 175 -58 209 58
<< nsubdiff >>
rect -323 219 -227 253
rect 227 219 323 253
rect -323 157 -289 219
rect 289 157 323 219
rect -323 -219 -289 -157
rect 289 -219 323 -157
rect -323 -253 -227 -219
rect 227 -253 323 -219
<< nsubdiffcont >>
rect -227 219 227 253
rect -323 -157 -289 157
rect 289 -157 323 157
rect -227 -253 227 -219
<< poly >>
rect -177 151 -111 167
rect -177 117 -161 151
rect -127 117 -111 151
rect -177 101 -111 117
rect 111 151 177 167
rect 111 117 127 151
rect 161 117 177 151
rect 111 101 177 117
rect -159 70 -129 101
rect -63 70 -33 96
rect 33 70 63 96
rect 129 70 159 101
rect -159 -96 -129 -70
rect -63 -101 -33 -70
rect 33 -101 63 -70
rect 129 -96 159 -70
rect -81 -117 81 -101
rect -81 -151 -65 -117
rect -31 -151 31 -117
rect 65 -151 81 -117
rect -81 -167 81 -151
<< polycont >>
rect -161 117 -127 151
rect 127 117 161 151
rect -65 -151 -31 -117
rect 31 -151 65 -117
<< locali >>
rect -323 219 -227 253
rect 227 219 323 253
rect -323 157 -289 219
rect 289 157 323 219
rect -177 117 -161 151
rect -127 117 -111 151
rect 111 117 127 151
rect 161 117 177 151
rect -209 58 -175 74
rect -209 -74 -175 -58
rect -113 58 -79 74
rect -113 -74 -79 -58
rect -17 58 17 74
rect -17 -74 17 -58
rect 79 58 113 74
rect 79 -74 113 -58
rect 175 58 209 74
rect 175 -74 209 -58
rect -81 -151 -65 -117
rect -31 -151 31 -117
rect 65 -151 81 -117
rect -323 -219 -289 -157
rect 289 -219 323 -157
rect -323 -253 -227 -219
rect 227 -253 323 -219
<< viali >>
rect -161 117 -127 151
rect 127 117 161 151
rect -209 -58 -175 58
rect -113 -58 -79 58
rect -17 -58 17 58
rect 79 -58 113 58
rect 175 -58 209 58
rect -65 -151 -31 -117
rect 31 -151 65 -117
<< metal1 >>
rect -173 151 -115 157
rect 115 151 173 157
rect -359 117 -161 151
rect -127 117 127 151
rect 161 117 359 151
rect -173 111 -115 117
rect 115 111 173 117
rect -225 58 -159 70
rect -225 -58 -218 58
rect -166 -58 -159 58
rect -225 -70 -159 -58
rect -129 58 -63 70
rect -129 -58 -122 58
rect -70 -58 -63 58
rect -129 -70 -63 -58
rect -33 58 33 70
rect -33 -58 -26 58
rect 26 -58 33 58
rect -33 -70 33 -58
rect 63 58 129 70
rect 63 -58 70 58
rect 122 -58 129 58
rect 63 -70 129 -58
rect 159 58 225 70
rect 159 -58 166 58
rect 218 -58 225 58
rect 159 -70 225 -58
rect -77 -117 77 -111
rect -77 -151 -65 -117
rect -31 -151 31 -117
rect 65 -151 359 -117
rect -77 -157 77 -151
rect -65 -289 -31 -157
<< via1 >>
rect -218 -58 -209 58
rect -209 -58 -175 58
rect -175 -58 -166 58
rect -122 -58 -113 58
rect -113 -58 -79 58
rect -79 -58 -70 58
rect -26 -58 -17 58
rect -17 -58 17 58
rect 17 -58 26 58
rect 70 -58 79 58
rect 79 -58 113 58
rect 113 -58 122 58
rect 166 -58 175 58
rect 175 -58 209 58
rect 209 -58 218 58
<< metal2 >>
rect -225 58 -159 70
rect -225 -58 -220 58
rect -164 -58 -159 58
rect -225 -70 -159 -58
rect -129 58 -63 70
rect -129 -58 -124 58
rect -68 -58 -63 58
rect -129 -70 -63 -58
rect -33 58 33 70
rect -33 -58 -26 58
rect 26 -58 33 58
rect -33 -70 33 -58
rect 63 58 129 70
rect 63 -58 68 58
rect 124 -58 129 58
rect 63 -70 129 -58
rect 159 58 225 70
rect 159 -58 164 58
rect 220 -58 225 58
rect 159 -70 225 -58
rect -17 -289 17 -70
<< via2 >>
rect -220 -58 -218 58
rect -218 -58 -166 58
rect -166 -58 -164 58
rect -124 -58 -122 58
rect -122 -58 -70 58
rect -70 -58 -68 58
rect 68 -58 70 58
rect 70 -58 122 58
rect 122 -58 124 58
rect 164 -58 166 58
rect 166 -58 218 58
rect 218 -58 220 58
<< metal3 >>
rect -359 58 359 70
rect -359 10 -220 58
rect -225 -58 -220 10
rect -164 -58 -124 58
rect -68 10 68 58
rect -68 -58 -63 10
rect -225 -70 -63 -58
rect 63 -58 68 10
rect 124 -58 164 58
rect 220 10 359 58
rect 220 -58 225 10
rect 63 -70 225 -58
<< properties >>
string FIXED_BBOX -306 -236 306 236
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.7 l 0.15 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
