magic
tech sky130A
timestamp 1668357910
<< metal3 >>
rect -425 -400 375 400
<< mimcap >>
rect -375 330 325 350
rect -375 -330 -355 330
rect 305 -330 325 330
rect -375 -350 325 -330
<< mimcapcontact >>
rect -355 -330 305 330
<< metal4 >>
rect -375 330 325 350
rect -375 -330 -355 330
rect 305 -330 325 330
rect -375 -350 325 -330
<< properties >>
string FIXED_BBOX -425 -400 375 400
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 7 l 7 val 103.32 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
