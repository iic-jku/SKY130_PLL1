magic
tech sky130A
magscale 1 2
timestamp 1666524377
<< error_s >>
rect 2870 1578 2928 1584
rect 2870 1544 2882 1578
rect 2870 1538 2928 1544
rect 1238 1310 1296 1316
rect 1238 1276 1250 1310
rect 1238 1270 1296 1276
<< metal1 >>
rect 2018 967 2390 1001
rect -42 539 0 581
rect 2172 534 2178 586
rect 2230 534 2236 586
rect 1826 138 2486 172
<< via1 >>
rect 2178 534 2230 586
<< metal2 >>
rect 26 1980 192 2050
rect 26 280 96 1980
rect 982 1427 1190 1497
rect 2976 1427 3184 1497
rect 982 919 1052 1427
rect 2528 918 2598 1329
rect 2178 586 2230 592
rect 3114 539 3156 581
rect 2178 528 2230 534
rect 3362 280 3432 1980
rect 26 210 234 280
rect 1875 210 2438 280
rect 2880 210 3716 280
use buffer  buffer_0 /foss/designs/ma2022
timestamp 1666523630
transform 1 0 0 0 1 0
box 0 0 2204 1138
use simple_inv  simple_inv_0 /foss/designs/ma2022
timestamp 1666523630
transform 1 0 2257 0 1 613
box -53 -613 857 525
use slope_p  sky130_fd_pr__pfet_01v8_BDAFKN_0 /foss/designs/ma2022
timestamp 1666523630
transform 1 0 2083 0 1 1427
box -1031 -289 1031 289
use tgate_1  tgate_1_0 /foss/designs/ma2022
timestamp 1666523630
transform 0 1 868 -1 0 2689
box -261 -952 919 1138
use tgate_1  tgate_1_1
timestamp 1666523630
transform 0 -1 3144 -1 0 2689
box -261 -952 919 1138
use tgate_1  tgate_1_2
timestamp 1666523630
transform -1 0 4425 0 1 632
box -261 -952 919 1138
<< labels >>
rlabel metal2 3114 539 3156 581 1 clk_out
rlabel metal1 -42 539 0 581 0 clk_in
<< end >>
