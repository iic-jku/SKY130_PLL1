magic
tech sky130A
magscale 1 2
timestamp 1668153059
<< metal1 >>
rect 1830 2866 1872 2908
rect 2140 2866 2182 2908
rect -866 1980 -858 2050
rect -788 1980 -621 2050
rect -551 1980 38 2050
rect 1402 1817 1454 1823
rect 1402 1759 1454 1765
rect 2558 1817 2610 1823
rect 2558 1759 2610 1765
rect 1407 1584 1449 1759
rect 2563 1584 2605 1759
rect 4602 1594 4644 1636
rect 1330 1538 2068 1584
rect 2482 1538 2644 1584
rect 3143 1427 3149 1497
rect 3219 1427 3503 1497
rect 3573 1427 3579 1497
rect 4504 1339 4574 1345
rect 3386 1316 3392 1319
rect 2097 1269 2508 1316
rect 2674 1270 3392 1316
rect 2466 1213 2508 1269
rect 3386 1267 3392 1270
rect 3444 1267 3450 1319
rect 3495 1213 3501 1218
rect 2466 1171 3501 1213
rect 3495 1166 3501 1171
rect 3553 1166 3559 1218
rect 3392 1118 3444 1124
rect 3392 1060 3444 1066
rect 4504 1118 4574 1269
rect 2657 588 2713 698
rect -625 539 -583 581
rect 1383 534 1389 586
rect 1441 534 1447 586
rect 2291 532 2297 588
rect 2353 532 2713 588
rect 2657 422 2713 532
rect 3114 441 3174 447
rect 3114 -240 3174 381
rect 3078 -259 3209 -240
rect 3078 -620 3099 -259
rect 3191 -620 3209 -259
rect 3395 -273 3441 1060
rect 4504 1042 4574 1048
rect 3386 -325 3392 -273
rect 3444 -325 3450 -273
rect 3078 -640 3209 -620
<< via1 >>
rect -858 1980 -788 2050
rect -621 1980 -551 2050
rect 1402 1765 1454 1817
rect 2558 1765 2610 1817
rect 3149 1427 3219 1497
rect 3503 1427 3573 1497
rect 3392 1267 3444 1319
rect 4504 1269 4574 1339
rect 3501 1166 3553 1218
rect 3392 1066 3444 1118
rect 1389 534 1441 586
rect 2297 532 2353 588
rect 3114 381 3174 441
rect 3099 -620 3191 -259
rect 4504 1048 4574 1118
rect 3392 -325 3444 -273
<< metal2 >>
rect 1407 2908 4686 2950
rect -737 2619 96 2689
rect 3916 2619 4166 2689
rect -858 2050 -788 2056
rect -858 280 -788 1980
rect -737 919 -667 2619
rect -621 2050 -551 2056
rect -625 1980 -621 2050
rect -551 1980 192 2050
rect 3214 1980 3381 2050
rect -621 1974 -551 1980
rect 1396 1765 1402 1817
rect 1454 1765 1460 1817
rect 2552 1765 2558 1817
rect 2610 1765 2616 1817
rect 3149 1497 3219 1503
rect 982 1427 1190 1497
rect 2976 1427 3149 1497
rect 3219 1427 3221 1497
rect 982 919 1052 1427
rect 3149 1421 3219 1427
rect 2652 919 2718 1329
rect -737 849 -650 919
rect 1279 849 1553 919
rect 1389 586 1441 592
rect 1389 528 1441 534
rect 2297 588 2353 594
rect 2297 526 2353 532
rect 2656 584 2714 779
rect 2656 536 3174 584
rect 2656 350 2714 536
rect 3114 441 3174 536
rect 3108 381 3114 441
rect 3174 381 3180 441
rect 3249 280 3319 1980
rect 4096 1806 4166 2619
rect 3637 1736 4574 1806
rect 3503 1497 3573 1503
rect 3637 1497 3707 1736
rect 3573 1427 3707 1497
rect 3503 1421 3573 1427
rect 4504 1339 4574 1736
rect 3392 1319 3444 1325
rect 4498 1269 4504 1339
rect 4574 1269 4580 1339
rect 3392 1261 3444 1267
rect 3395 1118 3441 1261
rect 3501 1218 3553 1224
rect 3501 1160 3553 1166
rect 4504 1118 4574 1120
rect 3386 1066 3392 1118
rect 3444 1066 3450 1118
rect 4498 1048 4504 1118
rect 4574 1048 4580 1118
rect 4504 632 4574 1048
rect 4355 562 4574 632
rect 4355 492 4425 562
rect -858 210 -554 280
rect 1087 210 1649 280
rect 2091 210 2466 280
rect 2903 210 3716 280
rect -858 -152 -788 210
rect -858 -252 1106 -152
rect 1206 -252 1215 -152
rect 3078 -259 3209 -240
rect 3078 -620 3099 -259
rect 3191 -620 3209 -259
rect 3392 -273 3444 -267
rect 4644 -278 4686 2908
rect 3444 -320 4686 -278
rect 3392 -331 3444 -325
rect 3078 -640 3209 -620
<< via2 >>
rect 1106 -252 1206 -152
rect 3099 -620 3191 -259
<< metal3 >>
rect 1101 -152 1211 -147
rect 1101 -252 1106 -152
rect 1206 -252 1211 -152
rect 1101 -257 1211 -252
rect 3078 -259 3209 -240
rect 3078 -620 3099 -259
rect 3191 -620 3209 -259
rect 3078 -640 3209 -620
<< via3 >>
rect 3099 -620 3191 -259
<< metal4 >>
rect 2706 -259 3209 -240
rect 2706 -620 3099 -259
rect 3191 -620 3209 -259
rect 2706 -640 3209 -620
use cap100f  cap100f_0
timestamp 1668153059
transform 1 0 2056 0 -1 -940
box -850 -800 750 800
use inv_buffer2  inv_buffer2_0
timestamp 1668153059
transform 1 0 -788 0 1 0
box 0 0 2204 1138
use inv_simple1  inv_simple1_0
timestamp 1668153059
transform 1 0 1468 0 1 613
box -53 -613 858 525
use sinv_n  sinv_n_0
timestamp 1668153059
transform 1 0 2685 0 1 280
box -359 -280 359 280
use slope_p  sky130_fd_pr__pfet_01v8_BDAFKN_0
timestamp 1668153059
transform 1 0 2083 0 1 1427
box -1031 -289 1031 289
use sinv_p2  sky130_fd_pr__pfet_01v8_X679XQ_0
timestamp 1668153059
transform 1 0 2685 0 1 849
box -359 -289 359 289
use tgate_1  tgate_1_0
timestamp 1668153059
transform 0 1 868 -1 0 2689
box -261 -952 919 1138
use tgate_1  tgate_1_1
timestamp 1668153059
transform 0 -1 3144 -1 0 2689
box -261 -952 919 1138
use tgate_1  tgate_1_2
timestamp 1668153059
transform -1 0 4425 0 1 632
box -261 -952 919 1138
<< labels >>
rlabel metal2 3114 539 3156 581 1 clk_out
port 1 n
rlabel metal1 4602 1594 4644 1636 3 bit1
port 2 n
rlabel metal1 2140 2866 2182 2908 7 bit0
port 3 n
rlabel metal1 1830 2866 1872 2908 3 bit2
port 4 n
rlabel metal1 3395 -261 3441 -215 0 vbias
port 5 n
rlabel metal1 -625 539 -583 581 0 clk_in
port 8 n
rlabel metal2 -737 1019 -667 1089 7 vdd
port 9 n
rlabel metal2 -858 1019 -788 1089 6 vss
port 10 n
<< end >>
