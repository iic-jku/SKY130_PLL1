magic
tech sky130A
magscale 1 2
timestamp 1668240031
<< viali >>
rect 1777 38505 1811 38539
rect 4721 38505 4755 38539
rect 7665 38505 7699 38539
rect 9873 38505 9907 38539
rect 11161 38505 11195 38539
rect 16313 38505 16347 38539
rect 22385 38505 22419 38539
rect 25881 38505 25915 38539
rect 27721 38505 27755 38539
rect 29929 38505 29963 38539
rect 34161 38505 34195 38539
rect 36921 38505 36955 38539
rect 12909 38437 12943 38471
rect 15301 38437 15335 38471
rect 30573 38437 30607 38471
rect 18429 38369 18463 38403
rect 19993 38369 20027 38403
rect 20729 38369 20763 38403
rect 1961 38301 1995 38335
rect 4905 38301 4939 38335
rect 7849 38301 7883 38335
rect 9689 38301 9723 38335
rect 10333 38301 10367 38335
rect 10977 38301 11011 38335
rect 12265 38301 12299 38335
rect 13093 38301 13127 38335
rect 13553 38301 13587 38335
rect 14657 38301 14691 38335
rect 15117 38301 15151 38335
rect 16129 38301 16163 38335
rect 17325 38301 17359 38335
rect 21005 38301 21039 38335
rect 22569 38301 22603 38335
rect 23029 38301 23063 38335
rect 23673 38301 23707 38335
rect 24777 38301 24811 38335
rect 25421 38301 25455 38335
rect 27997 38301 28031 38335
rect 28825 38301 28859 38335
rect 31217 38301 31251 38335
rect 31401 38301 31435 38335
rect 32505 38301 32539 38335
rect 32965 38301 32999 38335
rect 36737 38301 36771 38335
rect 13645 38233 13679 38267
rect 18245 38233 18279 38267
rect 19809 38233 19843 38267
rect 20913 38233 20947 38267
rect 29745 38233 29779 38267
rect 10517 38165 10551 38199
rect 12357 38165 12391 38199
rect 14473 38165 14507 38199
rect 17141 38165 17175 38199
rect 17785 38165 17819 38199
rect 18153 38165 18187 38199
rect 19441 38165 19475 38199
rect 19901 38165 19935 38199
rect 21373 38165 21407 38199
rect 23121 38165 23155 38199
rect 23765 38165 23799 38199
rect 24593 38165 24627 38199
rect 25237 38165 25271 38199
rect 27537 38165 27571 38199
rect 28733 38165 28767 38199
rect 29945 38165 29979 38199
rect 30113 38165 30147 38199
rect 31309 38165 31343 38199
rect 32413 38165 32447 38199
rect 33057 38165 33091 38199
rect 1593 37961 1627 37995
rect 5089 37961 5123 37995
rect 8125 37961 8159 37995
rect 10149 37961 10183 37995
rect 12449 37961 12483 37995
rect 13921 37961 13955 37995
rect 15761 37961 15795 37995
rect 18613 37961 18647 37995
rect 19257 37961 19291 37995
rect 21097 37961 21131 37995
rect 30021 37961 30055 37995
rect 34713 37961 34747 37995
rect 17141 37893 17175 37927
rect 20085 37893 20119 37927
rect 22293 37893 22327 37927
rect 24501 37893 24535 37927
rect 31493 37893 31527 37927
rect 1777 37825 1811 37859
rect 5273 37825 5307 37859
rect 8309 37825 8343 37859
rect 9597 37825 9631 37859
rect 10333 37825 10367 37859
rect 10793 37825 10827 37859
rect 11805 37825 11839 37859
rect 12817 37825 12851 37859
rect 12909 37825 12943 37859
rect 14289 37825 14323 37859
rect 15577 37825 15611 37859
rect 19073 37825 19107 37859
rect 20913 37825 20947 37859
rect 24225 37825 24259 37859
rect 26433 37825 26467 37859
rect 27261 37825 27295 37859
rect 28181 37825 28215 37859
rect 29561 37825 29595 37859
rect 34529 37825 34563 37859
rect 13093 37757 13127 37791
rect 14381 37757 14415 37791
rect 14473 37757 14507 37791
rect 16865 37757 16899 37791
rect 20177 37757 20211 37791
rect 20361 37757 20395 37791
rect 22017 37757 22051 37791
rect 23765 37757 23799 37791
rect 31769 37757 31803 37791
rect 33793 37757 33827 37791
rect 34069 37757 34103 37791
rect 11989 37689 12023 37723
rect 9413 37621 9447 37655
rect 10977 37621 11011 37655
rect 19717 37621 19751 37655
rect 25973 37621 26007 37655
rect 26525 37621 26559 37655
rect 27537 37621 27571 37655
rect 27721 37621 27755 37655
rect 28273 37621 28307 37655
rect 28641 37621 28675 37655
rect 29101 37621 29135 37655
rect 29469 37621 29503 37655
rect 32321 37621 32355 37655
rect 13461 37417 13495 37451
rect 14565 37417 14599 37451
rect 24041 37417 24075 37451
rect 28273 37417 28307 37451
rect 30205 37417 30239 37451
rect 27721 37349 27755 37383
rect 9413 37281 9447 37315
rect 15117 37281 15151 37315
rect 18337 37281 18371 37315
rect 23489 37281 23523 37315
rect 24961 37281 24995 37315
rect 25237 37281 25271 37315
rect 30021 37281 30055 37315
rect 8401 37213 8435 37247
rect 9137 37213 9171 37247
rect 11713 37213 11747 37247
rect 14933 37213 14967 37247
rect 15761 37213 15795 37247
rect 18521 37213 18555 37247
rect 19625 37213 19659 37247
rect 20269 37213 20303 37247
rect 22753 37213 22787 37247
rect 27905 37213 27939 37247
rect 28733 37213 28767 37247
rect 29193 37213 29227 37247
rect 29929 37213 29963 37247
rect 31033 37213 31067 37247
rect 33425 37213 33459 37247
rect 33517 37213 33551 37247
rect 11989 37145 12023 37179
rect 16037 37145 16071 37179
rect 18429 37145 18463 37179
rect 20545 37145 20579 37179
rect 23581 37145 23615 37179
rect 27997 37145 28031 37179
rect 28089 37145 28123 37179
rect 31309 37145 31343 37179
rect 8493 37077 8527 37111
rect 10885 37077 10919 37111
rect 15025 37077 15059 37111
rect 17509 37077 17543 37111
rect 18889 37077 18923 37111
rect 19809 37077 19843 37111
rect 22017 37077 22051 37111
rect 22569 37077 22603 37111
rect 23673 37077 23707 37111
rect 26709 37077 26743 37111
rect 28825 37077 28859 37111
rect 28917 37077 28951 37111
rect 32781 37077 32815 37111
rect 9781 36873 9815 36907
rect 11161 36873 11195 36907
rect 12633 36873 12667 36907
rect 13001 36873 13035 36907
rect 15577 36873 15611 36907
rect 16129 36873 16163 36907
rect 16957 36873 16991 36907
rect 17325 36873 17359 36907
rect 18153 36873 18187 36907
rect 20361 36873 20395 36907
rect 21373 36873 21407 36907
rect 24317 36873 24351 36907
rect 29015 36873 29049 36907
rect 10149 36805 10183 36839
rect 14105 36805 14139 36839
rect 19625 36805 19659 36839
rect 22385 36805 22419 36839
rect 24777 36805 24811 36839
rect 25881 36805 25915 36839
rect 27997 36805 28031 36839
rect 28917 36805 28951 36839
rect 29101 36805 29135 36839
rect 34069 36805 34103 36839
rect 9229 36737 9263 36771
rect 10977 36737 11011 36771
rect 12081 36737 12115 36771
rect 16313 36737 16347 36771
rect 17417 36737 17451 36771
rect 20545 36737 20579 36771
rect 21281 36737 21315 36771
rect 24685 36737 24719 36771
rect 25973 36737 26007 36771
rect 27169 36737 27203 36771
rect 29193 36737 29227 36771
rect 29837 36737 29871 36771
rect 30849 36737 30883 36771
rect 32321 36737 32355 36771
rect 10241 36669 10275 36703
rect 10425 36669 10459 36703
rect 13093 36669 13127 36703
rect 13277 36669 13311 36703
rect 13829 36669 13863 36703
rect 17509 36669 17543 36703
rect 19901 36669 19935 36703
rect 22109 36669 22143 36703
rect 24869 36669 24903 36703
rect 26065 36669 26099 36703
rect 29929 36669 29963 36703
rect 30205 36669 30239 36703
rect 25513 36601 25547 36635
rect 28365 36601 28399 36635
rect 9137 36533 9171 36567
rect 11989 36533 12023 36567
rect 23857 36533 23891 36567
rect 27261 36533 27295 36567
rect 28457 36533 28491 36567
rect 30757 36533 30791 36567
rect 9597 36329 9631 36363
rect 16957 36329 16991 36363
rect 18153 36329 18187 36363
rect 21925 36329 21959 36363
rect 23029 36329 23063 36363
rect 30113 36329 30147 36363
rect 33057 36329 33091 36363
rect 17601 36261 17635 36295
rect 25329 36261 25363 36295
rect 27997 36261 28031 36295
rect 28733 36261 28767 36295
rect 8493 36193 8527 36227
rect 10241 36193 10275 36227
rect 13461 36193 13495 36227
rect 13645 36193 13679 36227
rect 14933 36193 14967 36227
rect 18797 36193 18831 36227
rect 19901 36193 19935 36227
rect 23489 36193 23523 36227
rect 23581 36193 23615 36227
rect 24777 36193 24811 36227
rect 31309 36193 31343 36227
rect 7205 36125 7239 36159
rect 9965 36125 9999 36159
rect 10793 36125 10827 36159
rect 15209 36125 15243 36159
rect 17049 36125 17083 36159
rect 17693 36125 17727 36159
rect 18521 36125 18555 36159
rect 18613 36125 18647 36159
rect 20085 36125 20119 36159
rect 21833 36125 21867 36159
rect 24869 36125 24903 36159
rect 25973 36125 26007 36159
rect 26433 36125 26467 36159
rect 30205 36125 30239 36159
rect 30665 36125 30699 36159
rect 30849 36125 30883 36159
rect 33701 36125 33735 36159
rect 11069 36057 11103 36091
rect 13369 36057 13403 36091
rect 15117 36057 15151 36091
rect 27629 36057 27663 36091
rect 29009 36057 29043 36091
rect 31585 36057 31619 36091
rect 7297 35989 7331 36023
rect 7849 35989 7883 36023
rect 8217 35989 8251 36023
rect 8309 35989 8343 36023
rect 10057 35989 10091 36023
rect 12541 35989 12575 36023
rect 13001 35989 13035 36023
rect 15577 35989 15611 36023
rect 19993 35989 20027 36023
rect 20453 35989 20487 36023
rect 23397 35989 23431 36023
rect 24961 35989 24995 36023
rect 25789 35989 25823 36023
rect 26525 35989 26559 36023
rect 28089 35989 28123 36023
rect 28549 35989 28583 36023
rect 29745 35989 29779 36023
rect 30757 35989 30791 36023
rect 33609 35989 33643 36023
rect 10701 35785 10735 35819
rect 11161 35785 11195 35819
rect 13277 35785 13311 35819
rect 13645 35785 13679 35819
rect 15301 35785 15335 35819
rect 19165 35785 19199 35819
rect 20177 35785 20211 35819
rect 23489 35785 23523 35819
rect 23949 35785 23983 35819
rect 26617 35785 26651 35819
rect 27997 35785 28031 35819
rect 34069 35785 34103 35819
rect 12173 35717 12207 35751
rect 20085 35717 20119 35751
rect 23857 35717 23891 35751
rect 25145 35717 25179 35751
rect 28825 35717 28859 35751
rect 29837 35717 29871 35751
rect 30053 35717 30087 35751
rect 31585 35717 31619 35751
rect 32597 35717 32631 35751
rect 6561 35649 6595 35683
rect 7205 35649 7239 35683
rect 7849 35649 7883 35683
rect 10793 35649 10827 35683
rect 12081 35649 12115 35683
rect 14289 35649 14323 35683
rect 15393 35649 15427 35683
rect 16313 35649 16347 35683
rect 17877 35649 17911 35683
rect 19257 35649 19291 35683
rect 21189 35649 21223 35683
rect 22201 35649 22235 35683
rect 22937 35649 22971 35683
rect 24869 35649 24903 35683
rect 28089 35649 28123 35683
rect 28181 35649 28215 35683
rect 30849 35649 30883 35683
rect 31493 35649 31527 35683
rect 31677 35649 31711 35683
rect 32321 35649 32355 35683
rect 8125 35581 8159 35615
rect 10609 35581 10643 35615
rect 12265 35581 12299 35615
rect 13001 35581 13035 35615
rect 13185 35581 13219 35615
rect 15485 35581 15519 35615
rect 17969 35581 18003 35615
rect 18153 35581 18187 35615
rect 19901 35581 19935 35615
rect 24041 35581 24075 35615
rect 27721 35581 27755 35615
rect 27813 35581 27847 35615
rect 30665 35581 30699 35615
rect 7389 35513 7423 35547
rect 11713 35513 11747 35547
rect 14933 35513 14967 35547
rect 20545 35513 20579 35547
rect 29101 35513 29135 35547
rect 30205 35513 30239 35547
rect 6745 35445 6779 35479
rect 9597 35445 9631 35479
rect 14473 35445 14507 35479
rect 16129 35445 16163 35479
rect 17509 35445 17543 35479
rect 21005 35445 21039 35479
rect 22109 35445 22143 35479
rect 22753 35445 22787 35479
rect 28365 35445 28399 35479
rect 29285 35445 29319 35479
rect 30021 35445 30055 35479
rect 31033 35445 31067 35479
rect 6910 35241 6944 35275
rect 8401 35241 8435 35275
rect 10333 35241 10367 35275
rect 18245 35241 18279 35275
rect 22385 35241 22419 35275
rect 23305 35241 23339 35275
rect 27261 35241 27295 35275
rect 28181 35241 28215 35275
rect 28365 35241 28399 35275
rect 28641 35241 28675 35275
rect 29929 35241 29963 35275
rect 33517 35241 33551 35275
rect 6653 35105 6687 35139
rect 9597 35105 9631 35139
rect 9781 35105 9815 35139
rect 10977 35105 11011 35139
rect 14289 35105 14323 35139
rect 16497 35105 16531 35139
rect 19901 35105 19935 35139
rect 19993 35105 20027 35139
rect 20637 35105 20671 35139
rect 23857 35105 23891 35139
rect 24777 35105 24811 35139
rect 26341 35105 26375 35139
rect 28273 35105 28307 35139
rect 32965 35105 32999 35139
rect 1777 35037 1811 35071
rect 10793 35037 10827 35071
rect 11621 35037 11655 35071
rect 12265 35037 12299 35071
rect 12909 35037 12943 35071
rect 13553 35037 13587 35071
rect 18889 35037 18923 35071
rect 24961 35037 24995 35071
rect 26249 35037 26283 35071
rect 26985 35037 27019 35071
rect 27905 35037 27939 35071
rect 28089 35037 28123 35071
rect 30205 35037 30239 35071
rect 33609 35037 33643 35071
rect 36921 35037 36955 35071
rect 14565 34969 14599 35003
rect 16773 34969 16807 35003
rect 18797 34969 18831 35003
rect 20913 34969 20947 35003
rect 23673 34969 23707 35003
rect 26157 34969 26191 35003
rect 32689 34969 32723 35003
rect 1593 34901 1627 34935
rect 9137 34901 9171 34935
rect 9505 34901 9539 34935
rect 10701 34901 10735 34935
rect 11805 34901 11839 34935
rect 12357 34901 12391 34935
rect 13001 34901 13035 34935
rect 13737 34901 13771 34935
rect 16037 34901 16071 34935
rect 19441 34901 19475 34935
rect 19809 34901 19843 34935
rect 23765 34901 23799 34935
rect 24869 34901 24903 34935
rect 25329 34901 25363 34935
rect 25789 34901 25823 34935
rect 27445 34901 27479 34935
rect 29745 34901 29779 34935
rect 31217 34901 31251 34935
rect 37105 34901 37139 34935
rect 8493 34697 8527 34731
rect 8861 34697 8895 34731
rect 8953 34697 8987 34731
rect 11713 34697 11747 34731
rect 13001 34697 13035 34731
rect 15577 34697 15611 34731
rect 16313 34697 16347 34731
rect 18061 34697 18095 34731
rect 18521 34697 18555 34731
rect 23949 34697 23983 34731
rect 24777 34697 24811 34731
rect 24869 34697 24903 34731
rect 25697 34697 25731 34731
rect 28273 34697 28307 34731
rect 28641 34697 28675 34731
rect 30934 34697 30968 34731
rect 31585 34697 31619 34731
rect 22477 34629 22511 34663
rect 28181 34629 28215 34663
rect 31033 34629 31067 34663
rect 32321 34629 32355 34663
rect 10333 34561 10367 34595
rect 10977 34561 11011 34595
rect 12081 34561 12115 34595
rect 14749 34561 14783 34595
rect 15669 34561 15703 34595
rect 16129 34561 16163 34595
rect 17417 34561 17451 34595
rect 18429 34561 18463 34595
rect 19441 34561 19475 34595
rect 25605 34561 25639 34595
rect 26433 34561 26467 34595
rect 27905 34561 27939 34595
rect 28365 34561 28399 34595
rect 29285 34561 29319 34595
rect 29929 34561 29963 34595
rect 30757 34561 30791 34595
rect 30849 34561 30883 34595
rect 31493 34561 31527 34595
rect 31677 34561 31711 34595
rect 9137 34493 9171 34527
rect 11069 34493 11103 34527
rect 12173 34493 12207 34527
rect 12357 34493 12391 34527
rect 18613 34493 18647 34527
rect 21189 34493 21223 34527
rect 22201 34493 22235 34527
rect 24961 34493 24995 34527
rect 29193 34493 29227 34527
rect 30021 34493 30055 34527
rect 30297 34425 30331 34459
rect 33609 34425 33643 34459
rect 10517 34357 10551 34391
rect 14491 34357 14525 34391
rect 17509 34357 17543 34391
rect 19698 34357 19732 34391
rect 24409 34357 24443 34391
rect 26249 34357 26283 34391
rect 27997 34357 28031 34391
rect 12633 34153 12667 34187
rect 15025 34153 15059 34187
rect 18245 34153 18279 34187
rect 20821 34153 20855 34187
rect 26709 34153 26743 34187
rect 27813 34153 27847 34187
rect 33149 34153 33183 34187
rect 19533 34085 19567 34119
rect 8401 34017 8435 34051
rect 9597 34017 9631 34051
rect 9689 34017 9723 34051
rect 10701 34017 10735 34051
rect 13185 34017 13219 34051
rect 14381 34017 14415 34051
rect 16129 34017 16163 34051
rect 20085 34017 20119 34051
rect 23397 34017 23431 34051
rect 24961 34017 24995 34051
rect 25237 34017 25271 34051
rect 10425 33949 10459 33983
rect 13093 33949 13127 33983
rect 15945 33949 15979 33983
rect 16773 33949 16807 33983
rect 17417 33949 17451 33983
rect 18061 33949 18095 33983
rect 18705 33949 18739 33983
rect 20913 33949 20947 33983
rect 22201 33949 22235 33983
rect 23213 33949 23247 33983
rect 27997 33949 28031 33983
rect 28089 33949 28123 33983
rect 28273 33949 28307 33983
rect 28365 33949 28399 33983
rect 29929 33949 29963 33983
rect 32597 33949 32631 33983
rect 33241 33949 33275 33983
rect 14565 33881 14599 33915
rect 19993 33881 20027 33915
rect 32321 33881 32355 33915
rect 7849 33813 7883 33847
rect 8217 33813 8251 33847
rect 8309 33813 8343 33847
rect 9137 33813 9171 33847
rect 9505 33813 9539 33847
rect 12173 33813 12207 33847
rect 13001 33813 13035 33847
rect 14657 33813 14691 33847
rect 15577 33813 15611 33847
rect 16037 33813 16071 33847
rect 16865 33813 16899 33847
rect 17601 33813 17635 33847
rect 18889 33813 18923 33847
rect 19901 33813 19935 33847
rect 22293 33813 22327 33847
rect 22845 33813 22879 33847
rect 23305 33813 23339 33847
rect 29837 33813 29871 33847
rect 30849 33813 30883 33847
rect 9597 33609 9631 33643
rect 10793 33609 10827 33643
rect 15577 33609 15611 33643
rect 15945 33609 15979 33643
rect 19073 33609 19107 33643
rect 32413 33609 32447 33643
rect 33057 33609 33091 33643
rect 10425 33541 10459 33575
rect 12541 33541 12575 33575
rect 17601 33541 17635 33575
rect 19625 33541 19659 33575
rect 30665 33541 30699 33575
rect 7389 33473 7423 33507
rect 7849 33473 7883 33507
rect 10333 33473 10367 33507
rect 14933 33473 14967 33507
rect 20453 33473 20487 33507
rect 22017 33473 22051 33507
rect 24225 33473 24259 33507
rect 24869 33473 24903 33507
rect 29377 33473 29411 33507
rect 30573 33473 30607 33507
rect 30757 33473 30791 33507
rect 31217 33473 31251 33507
rect 31401 33473 31435 33507
rect 32321 33473 32355 33507
rect 32505 33473 32539 33507
rect 33149 33473 33183 33507
rect 8125 33405 8159 33439
rect 10241 33405 10275 33439
rect 12265 33405 12299 33439
rect 14013 33405 14047 33439
rect 16037 33405 16071 33439
rect 16221 33405 16255 33439
rect 17325 33405 17359 33439
rect 22293 33405 22327 33439
rect 25145 33405 25179 33439
rect 28089 33405 28123 33439
rect 28549 33405 28583 33439
rect 29193 33405 29227 33439
rect 31309 33405 31343 33439
rect 24409 33337 24443 33371
rect 28365 33337 28399 33371
rect 29009 33337 29043 33371
rect 29285 33337 29319 33371
rect 7205 33269 7239 33303
rect 15117 33269 15151 33303
rect 23765 33269 23799 33303
rect 26617 33269 26651 33303
rect 29193 33269 29227 33303
rect 8493 33065 8527 33099
rect 9597 33065 9631 33099
rect 12357 33065 12391 33099
rect 14657 33065 14691 33099
rect 16110 33065 16144 33099
rect 18153 33065 18187 33099
rect 24593 33065 24627 33099
rect 26065 33065 26099 33099
rect 26709 33065 26743 33099
rect 30481 33065 30515 33099
rect 34345 33065 34379 33099
rect 21189 32997 21223 33031
rect 27721 32997 27755 33031
rect 27905 32997 27939 33031
rect 31033 32997 31067 33031
rect 7021 32929 7055 32963
rect 10057 32929 10091 32963
rect 10241 32929 10275 32963
rect 11713 32929 11747 32963
rect 11897 32929 11931 32963
rect 15209 32929 15243 32963
rect 15853 32929 15887 32963
rect 18613 32929 18647 32963
rect 18705 32929 18739 32963
rect 19441 32929 19475 32963
rect 22569 32929 22603 32963
rect 23765 32929 23799 32963
rect 25145 32929 25179 32963
rect 27445 32929 27479 32963
rect 28457 32929 28491 32963
rect 28549 32929 28583 32963
rect 30113 32929 30147 32963
rect 33701 32929 33735 32963
rect 6745 32861 6779 32895
rect 10977 32861 11011 32895
rect 13277 32861 13311 32895
rect 15025 32861 15059 32895
rect 21833 32861 21867 32895
rect 23581 32861 23615 32895
rect 25053 32861 25087 32895
rect 26157 32861 26191 32895
rect 26801 32861 26835 32895
rect 28641 32861 28675 32895
rect 28733 32861 28767 32895
rect 30297 32861 30331 32895
rect 32781 32861 32815 32895
rect 9965 32793 9999 32827
rect 19717 32793 19751 32827
rect 23673 32793 23707 32827
rect 32505 32793 32539 32827
rect 33977 32793 34011 32827
rect 11069 32725 11103 32759
rect 11989 32725 12023 32759
rect 13185 32725 13219 32759
rect 15117 32725 15151 32759
rect 17601 32725 17635 32759
rect 18521 32725 18555 32759
rect 23213 32725 23247 32759
rect 24961 32725 24995 32759
rect 28917 32725 28951 32759
rect 33885 32725 33919 32759
rect 7389 32521 7423 32555
rect 14105 32521 14139 32555
rect 19165 32521 19199 32555
rect 19625 32521 19659 32555
rect 20453 32521 20487 32555
rect 22661 32521 22695 32555
rect 23673 32521 23707 32555
rect 24777 32521 24811 32555
rect 25237 32521 25271 32555
rect 30113 32521 30147 32555
rect 31217 32521 31251 32555
rect 33057 32521 33091 32555
rect 7941 32453 7975 32487
rect 27813 32453 27847 32487
rect 29653 32453 29687 32487
rect 34345 32453 34379 32487
rect 6561 32385 6595 32419
rect 7205 32385 7239 32419
rect 8033 32385 8067 32419
rect 8493 32385 8527 32419
rect 9321 32385 9355 32419
rect 10333 32385 10367 32419
rect 10977 32385 11011 32419
rect 12081 32385 12115 32419
rect 13369 32385 13403 32419
rect 17049 32385 17083 32419
rect 18061 32385 18095 32419
rect 19533 32385 19567 32419
rect 20361 32385 20395 32419
rect 21281 32385 21315 32419
rect 22201 32385 22235 32419
rect 22845 32385 22879 32419
rect 24869 32385 24903 32419
rect 25881 32385 25915 32419
rect 26525 32385 26559 32419
rect 27353 32385 27387 32419
rect 29929 32385 29963 32419
rect 31125 32385 31159 32419
rect 31401 32385 31435 32419
rect 32505 32385 32539 32419
rect 32965 32385 32999 32419
rect 33149 32385 33183 32419
rect 33793 32385 33827 32419
rect 34253 32385 34287 32419
rect 12173 32317 12207 32351
rect 12265 32317 12299 32351
rect 13461 32317 13495 32351
rect 15853 32317 15887 32351
rect 19717 32317 19751 32351
rect 23765 32317 23799 32351
rect 23949 32317 23983 32351
rect 24685 32317 24719 32351
rect 28273 32317 28307 32351
rect 28733 32317 28767 32351
rect 29193 32317 29227 32351
rect 29745 32317 29779 32351
rect 28181 32249 28215 32283
rect 29009 32249 29043 32283
rect 31401 32249 31435 32283
rect 32413 32249 32447 32283
rect 6745 32181 6779 32215
rect 8677 32181 8711 32215
rect 9229 32181 9263 32215
rect 10425 32181 10459 32215
rect 11161 32181 11195 32215
rect 11713 32181 11747 32215
rect 15589 32181 15623 32215
rect 16865 32181 16899 32215
rect 18153 32181 18187 32215
rect 21373 32181 21407 32215
rect 22017 32181 22051 32215
rect 23305 32181 23339 32215
rect 25697 32181 25731 32215
rect 26433 32181 26467 32215
rect 27261 32181 27295 32215
rect 29929 32181 29963 32215
rect 33701 32181 33735 32215
rect 7297 31977 7331 32011
rect 7849 31977 7883 32011
rect 9321 31977 9355 32011
rect 12246 31977 12280 32011
rect 13737 31977 13771 32011
rect 15025 31977 15059 32011
rect 20992 31977 21026 32011
rect 22937 31977 22971 32011
rect 27813 31977 27847 32011
rect 33057 31977 33091 32011
rect 11529 31909 11563 31943
rect 22477 31909 22511 31943
rect 8401 31841 8435 31875
rect 10057 31841 10091 31875
rect 11989 31841 12023 31875
rect 14381 31841 14415 31875
rect 14565 31841 14599 31875
rect 16129 31841 16163 31875
rect 18889 31841 18923 31875
rect 20729 31841 20763 31875
rect 23489 31841 23523 31875
rect 24961 31841 24995 31875
rect 26433 31841 26467 31875
rect 29193 31841 29227 31875
rect 31309 31841 31343 31875
rect 1777 31773 1811 31807
rect 6561 31773 6595 31807
rect 7205 31773 7239 31807
rect 9137 31773 9171 31807
rect 9781 31773 9815 31807
rect 17141 31773 17175 31807
rect 19625 31773 19659 31807
rect 20085 31773 20119 31807
rect 20177 31773 20211 31807
rect 23305 31773 23339 31807
rect 23397 31773 23431 31807
rect 24685 31773 24719 31807
rect 26985 31773 27019 31807
rect 27077 31773 27111 31807
rect 27629 31773 27663 31807
rect 28089 31773 28123 31807
rect 28549 31773 28583 31807
rect 28733 31773 28767 31807
rect 28825 31773 28859 31807
rect 28917 31773 28951 31807
rect 29837 31773 29871 31807
rect 29929 31773 29963 31807
rect 30021 31773 30055 31807
rect 30205 31773 30239 31807
rect 30849 31773 30883 31807
rect 33701 31773 33735 31807
rect 33793 31773 33827 31807
rect 36921 31773 36955 31807
rect 15945 31705 15979 31739
rect 17417 31705 17451 31739
rect 31585 31705 31619 31739
rect 1593 31637 1627 31671
rect 6653 31637 6687 31671
rect 8217 31637 8251 31671
rect 8309 31637 8343 31671
rect 14657 31637 14691 31671
rect 15577 31637 15611 31671
rect 16037 31637 16071 31671
rect 19441 31637 19475 31671
rect 27997 31637 28031 31671
rect 30757 31637 30791 31671
rect 37105 31637 37139 31671
rect 7205 31433 7239 31467
rect 10425 31433 10459 31467
rect 10793 31433 10827 31467
rect 11897 31433 11931 31467
rect 17049 31433 17083 31467
rect 17877 31433 17911 31467
rect 18705 31433 18739 31467
rect 19073 31433 19107 31467
rect 22845 31433 22879 31467
rect 24225 31433 24259 31467
rect 33793 31433 33827 31467
rect 34621 31433 34655 31467
rect 7941 31365 7975 31399
rect 10885 31365 10919 31399
rect 14289 31365 14323 31399
rect 24961 31365 24995 31399
rect 30389 31365 30423 31399
rect 31017 31365 31051 31399
rect 31217 31365 31251 31399
rect 32689 31365 32723 31399
rect 7021 31297 7055 31331
rect 11713 31297 11747 31331
rect 12357 31297 12391 31331
rect 16865 31297 16899 31331
rect 17969 31297 18003 31331
rect 20729 31297 20763 31331
rect 21281 31297 21315 31331
rect 22753 31297 22787 31331
rect 24041 31297 24075 31331
rect 27997 31297 28031 31331
rect 32597 31297 32631 31331
rect 33609 31297 33643 31331
rect 34437 31297 34471 31331
rect 7665 31229 7699 31263
rect 10977 31229 11011 31263
rect 13185 31229 13219 31263
rect 14013 31229 14047 31263
rect 18153 31229 18187 31263
rect 19165 31229 19199 31263
rect 19349 31229 19383 31263
rect 22661 31229 22695 31263
rect 24685 31229 24719 31263
rect 32413 31229 32447 31263
rect 17509 31161 17543 31195
rect 20453 31161 20487 31195
rect 26433 31161 26467 31195
rect 27537 31161 27571 31195
rect 30849 31161 30883 31195
rect 33057 31161 33091 31195
rect 9413 31093 9447 31127
rect 15761 31093 15795 31127
rect 21373 31093 21407 31127
rect 23213 31093 23247 31127
rect 27905 31093 27939 31127
rect 29101 31093 29135 31127
rect 31033 31093 31067 31127
rect 8217 30889 8251 30923
rect 11805 30889 11839 30923
rect 14749 30889 14783 30923
rect 15945 30889 15979 30923
rect 19441 30889 19475 30923
rect 21189 30889 21223 30923
rect 24593 30889 24627 30923
rect 28733 30889 28767 30923
rect 29745 30889 29779 30923
rect 30113 30889 30147 30923
rect 32689 30889 32723 30923
rect 34345 30889 34379 30923
rect 13369 30821 13403 30855
rect 28917 30821 28951 30855
rect 9965 30753 9999 30787
rect 12265 30753 12299 30787
rect 12357 30753 12391 30787
rect 15301 30753 15335 30787
rect 17417 30753 17451 30787
rect 18705 30753 18739 30787
rect 19901 30753 19935 30787
rect 19993 30753 20027 30787
rect 25145 30753 25179 30787
rect 30941 30753 30975 30787
rect 31217 30753 31251 30787
rect 33701 30753 33735 30787
rect 6469 30685 6503 30719
rect 9229 30685 9263 30719
rect 12173 30685 12207 30719
rect 15117 30685 15151 30719
rect 17693 30685 17727 30719
rect 18889 30685 18923 30719
rect 19809 30685 19843 30719
rect 22937 30685 22971 30719
rect 23581 30685 23615 30719
rect 24961 30685 24995 30719
rect 25973 30685 26007 30719
rect 26617 30685 26651 30719
rect 27353 30685 27387 30719
rect 27446 30685 27480 30719
rect 27629 30685 27663 30719
rect 27859 30685 27893 30719
rect 28457 30685 28491 30719
rect 30205 30685 30239 30719
rect 6745 30617 6779 30651
rect 10793 30617 10827 30651
rect 13645 30617 13679 30651
rect 15209 30617 15243 30651
rect 22661 30617 22695 30651
rect 25053 30617 25087 30651
rect 27721 30617 27755 30651
rect 9321 30549 9355 30583
rect 23397 30549 23431 30583
rect 25789 30549 25823 30583
rect 26525 30549 26559 30583
rect 27997 30549 28031 30583
rect 33885 30549 33919 30583
rect 33977 30549 34011 30583
rect 9597 30345 9631 30379
rect 25421 30345 25455 30379
rect 27261 30345 27295 30379
rect 7297 30277 7331 30311
rect 8493 30277 8527 30311
rect 9505 30277 9539 30311
rect 10793 30277 10827 30311
rect 13277 30277 13311 30311
rect 14841 30277 14875 30311
rect 16221 30277 16255 30311
rect 17233 30277 17267 30311
rect 17325 30277 17359 30311
rect 19349 30277 19383 30311
rect 22201 30277 22235 30311
rect 28733 30277 28767 30311
rect 29621 30277 29655 30311
rect 29837 30277 29871 30311
rect 7205 30209 7239 30243
rect 8401 30209 8435 30243
rect 10885 30209 10919 30243
rect 12357 30209 12391 30243
rect 13185 30209 13219 30243
rect 14473 30209 14507 30243
rect 15485 30209 15519 30243
rect 16313 30209 16347 30243
rect 18245 30209 18279 30243
rect 18521 30209 18555 30243
rect 19073 30209 19107 30243
rect 21465 30209 21499 30243
rect 22477 30209 22511 30243
rect 23857 30209 23891 30243
rect 23949 30209 23983 30243
rect 25053 30209 25087 30243
rect 26249 30209 26283 30243
rect 27537 30209 27571 30243
rect 27626 30209 27660 30243
rect 27726 30209 27760 30243
rect 27905 30209 27939 30243
rect 28544 30209 28578 30243
rect 28641 30209 28675 30243
rect 28861 30209 28895 30243
rect 29009 30209 29043 30243
rect 30665 30209 30699 30243
rect 31493 30209 31527 30243
rect 32321 30209 32355 30243
rect 33681 30209 33715 30243
rect 7481 30141 7515 30175
rect 8677 30141 8711 30175
rect 9413 30141 9447 30175
rect 10977 30141 11011 30175
rect 12173 30141 12207 30175
rect 13461 30141 13495 30175
rect 17417 30141 17451 30175
rect 20821 30141 20855 30175
rect 24041 30141 24075 30175
rect 24869 30141 24903 30175
rect 24961 30141 24995 30175
rect 30573 30141 30607 30175
rect 31033 30141 31067 30175
rect 32597 30141 32631 30175
rect 33425 30141 33459 30175
rect 6837 30073 6871 30107
rect 8033 30073 8067 30107
rect 10425 30073 10459 30107
rect 29469 30073 29503 30107
rect 34805 30073 34839 30107
rect 9965 30005 9999 30039
rect 12817 30005 12851 30039
rect 15301 30005 15335 30039
rect 16865 30005 16899 30039
rect 21281 30005 21315 30039
rect 23489 30005 23523 30039
rect 25973 30005 26007 30039
rect 28365 30005 28399 30039
rect 29653 30005 29687 30039
rect 31585 30005 31619 30039
rect 12909 29801 12943 29835
rect 14565 29801 14599 29835
rect 15761 29801 15795 29835
rect 19717 29801 19751 29835
rect 23121 29801 23155 29835
rect 26709 29801 26743 29835
rect 28457 29801 28491 29835
rect 30941 29801 30975 29835
rect 33057 29801 33091 29835
rect 7849 29733 7883 29767
rect 22661 29733 22695 29767
rect 8309 29665 8343 29699
rect 8401 29665 8435 29699
rect 10241 29665 10275 29699
rect 10425 29665 10459 29699
rect 11437 29665 11471 29699
rect 16405 29665 16439 29699
rect 18245 29665 18279 29699
rect 20913 29665 20947 29699
rect 23581 29665 23615 29699
rect 23673 29665 23707 29699
rect 25237 29665 25271 29699
rect 27997 29665 28031 29699
rect 28089 29665 28123 29699
rect 28917 29665 28951 29699
rect 33885 29665 33919 29699
rect 5917 29597 5951 29631
rect 6561 29597 6595 29631
rect 7205 29597 7239 29631
rect 9137 29597 9171 29631
rect 10149 29597 10183 29631
rect 11161 29597 11195 29631
rect 13737 29597 13771 29631
rect 17049 29597 17083 29631
rect 19809 29597 19843 29631
rect 23489 29597 23523 29631
rect 24961 29597 24995 29631
rect 27721 29597 27755 29631
rect 27905 29597 27939 29631
rect 28273 29597 28307 29631
rect 29101 29597 29135 29631
rect 29193 29597 29227 29631
rect 29745 29597 29779 29631
rect 30113 29597 30147 29631
rect 31769 29597 31803 29631
rect 32229 29597 32263 29631
rect 32873 29597 32907 29631
rect 33517 29597 33551 29631
rect 33701 29597 33735 29631
rect 9229 29529 9263 29563
rect 14657 29529 14691 29563
rect 17325 29529 17359 29563
rect 21189 29529 21223 29563
rect 28917 29529 28951 29563
rect 29929 29529 29963 29563
rect 30021 29529 30055 29563
rect 30757 29529 30791 29563
rect 31677 29529 31711 29563
rect 6101 29461 6135 29495
rect 6653 29461 6687 29495
rect 7389 29461 7423 29495
rect 8217 29461 8251 29495
rect 9781 29461 9815 29495
rect 13645 29461 13679 29495
rect 16129 29461 16163 29495
rect 16221 29461 16255 29495
rect 18429 29461 18463 29495
rect 18521 29461 18555 29495
rect 18889 29461 18923 29495
rect 30297 29461 30331 29495
rect 30957 29461 30991 29495
rect 31125 29461 31159 29495
rect 32413 29461 32447 29495
rect 11069 29257 11103 29291
rect 17233 29257 17267 29291
rect 21373 29257 21407 29291
rect 22753 29257 22787 29291
rect 23581 29257 23615 29291
rect 29101 29257 29135 29291
rect 29561 29257 29595 29291
rect 29745 29257 29779 29291
rect 31309 29257 31343 29291
rect 31769 29257 31803 29291
rect 33057 29257 33091 29291
rect 34897 29257 34931 29291
rect 6837 29189 6871 29223
rect 9597 29189 9631 29223
rect 19533 29189 19567 29223
rect 27537 29189 27571 29223
rect 31401 29189 31435 29223
rect 34192 29189 34226 29223
rect 6561 29121 6595 29155
rect 11897 29121 11931 29155
rect 19625 29121 19659 29155
rect 20269 29121 20303 29155
rect 21465 29121 21499 29155
rect 23949 29121 23983 29155
rect 27445 29121 27479 29155
rect 28365 29121 28399 29155
rect 28549 29121 28583 29155
rect 28917 29121 28951 29155
rect 29686 29121 29720 29155
rect 30113 29121 30147 29155
rect 30205 29121 30239 29155
rect 32321 29121 32355 29155
rect 35081 29121 35115 29155
rect 9321 29053 9355 29087
rect 12357 29053 12391 29087
rect 12633 29053 12667 29087
rect 14565 29053 14599 29087
rect 14841 29053 14875 29087
rect 18981 29053 19015 29087
rect 22845 29053 22879 29087
rect 23029 29053 23063 29087
rect 24041 29053 24075 29087
rect 24133 29053 24167 29087
rect 24869 29053 24903 29087
rect 25145 29053 25179 29087
rect 28641 29053 28675 29087
rect 28733 29053 28767 29087
rect 31125 29053 31159 29087
rect 34437 29053 34471 29087
rect 11805 28985 11839 29019
rect 20085 28985 20119 29019
rect 26617 28985 26651 29019
rect 8309 28917 8343 28951
rect 14105 28917 14139 28951
rect 16313 28917 16347 28951
rect 18723 28917 18757 28951
rect 22385 28917 22419 28951
rect 32505 28917 32539 28951
rect 10517 28713 10551 28747
rect 15577 28713 15611 28747
rect 16865 28713 16899 28747
rect 25789 28713 25823 28747
rect 26525 28713 26559 28747
rect 29009 28713 29043 28747
rect 30297 28713 30331 28747
rect 31125 28713 31159 28747
rect 33885 28713 33919 28747
rect 14289 28645 14323 28679
rect 25329 28645 25363 28679
rect 8401 28577 8435 28611
rect 9597 28577 9631 28611
rect 9689 28577 9723 28611
rect 11161 28577 11195 28611
rect 12817 28577 12851 28611
rect 14933 28577 14967 28611
rect 17509 28577 17543 28611
rect 18613 28577 18647 28611
rect 18705 28577 18739 28611
rect 20453 28577 20487 28611
rect 22201 28577 22235 28611
rect 23857 28577 23891 28611
rect 24777 28577 24811 28611
rect 28549 28577 28583 28611
rect 28641 28577 28675 28611
rect 33241 28577 33275 28611
rect 7205 28509 7239 28543
rect 10333 28509 10367 28543
rect 13737 28509 13771 28543
rect 15485 28509 15519 28543
rect 16313 28509 16347 28543
rect 17233 28509 17267 28543
rect 19993 28509 20027 28543
rect 23581 28509 23615 28543
rect 24869 28509 24903 28543
rect 25973 28509 26007 28543
rect 26617 28509 26651 28543
rect 28273 28509 28307 28543
rect 28457 28509 28491 28543
rect 28825 28509 28859 28543
rect 29745 28509 29779 28543
rect 29837 28509 29871 28543
rect 30021 28509 30055 28543
rect 30113 28509 30147 28543
rect 32505 28509 32539 28543
rect 33425 28509 33459 28543
rect 34897 28509 34931 28543
rect 35081 28509 35115 28543
rect 35725 28509 35759 28543
rect 8125 28441 8159 28475
rect 12541 28441 12575 28475
rect 20729 28441 20763 28475
rect 24961 28441 24995 28475
rect 32260 28441 32294 28475
rect 7021 28373 7055 28407
rect 7757 28373 7791 28407
rect 8217 28373 8251 28407
rect 9137 28373 9171 28407
rect 9505 28373 9539 28407
rect 11253 28373 11287 28407
rect 11345 28373 11379 28407
rect 11713 28373 11747 28407
rect 13553 28373 13587 28407
rect 14657 28373 14691 28407
rect 14749 28373 14783 28407
rect 16129 28373 16163 28407
rect 17325 28373 17359 28407
rect 18153 28373 18187 28407
rect 18521 28373 18555 28407
rect 19901 28373 19935 28407
rect 23213 28373 23247 28407
rect 23673 28373 23707 28407
rect 33517 28373 33551 28407
rect 34989 28373 35023 28407
rect 35541 28373 35575 28407
rect 8309 28169 8343 28203
rect 11161 28169 11195 28203
rect 12357 28169 12391 28203
rect 14197 28169 14231 28203
rect 15393 28169 15427 28203
rect 16865 28169 16899 28203
rect 18245 28169 18279 28203
rect 20913 28169 20947 28203
rect 28733 28169 28767 28203
rect 29837 28169 29871 28203
rect 34069 28169 34103 28203
rect 6837 28101 6871 28135
rect 8861 28101 8895 28135
rect 12725 28101 12759 28135
rect 15761 28101 15795 28135
rect 17325 28101 17359 28135
rect 18981 28101 19015 28135
rect 25329 28101 25363 28135
rect 32413 28101 32447 28135
rect 35173 28101 35207 28135
rect 1777 28033 1811 28067
rect 6561 28033 6595 28067
rect 8769 28033 8803 28067
rect 9413 28033 9447 28067
rect 11897 28033 11931 28067
rect 12817 28033 12851 28067
rect 13553 28033 13587 28067
rect 14565 28033 14599 28067
rect 14657 28033 14691 28067
rect 17233 28033 17267 28067
rect 18061 28033 18095 28067
rect 21097 28033 21131 28067
rect 22201 28033 22235 28067
rect 23029 28033 23063 28067
rect 24225 28033 24259 28067
rect 24317 28033 24351 28067
rect 25421 28033 25455 28067
rect 26433 28033 26467 28067
rect 27905 28033 27939 28067
rect 29009 28033 29043 28067
rect 29285 28033 29319 28067
rect 29745 28033 29779 28067
rect 30021 28033 30055 28067
rect 30205 28033 30239 28067
rect 30665 28033 30699 28067
rect 31033 28033 31067 28067
rect 31217 28033 31251 28067
rect 33425 28033 33459 28067
rect 33517 28033 33551 28067
rect 33977 28033 34011 28067
rect 34161 28033 34195 28067
rect 9689 27965 9723 27999
rect 12909 27965 12943 27999
rect 14841 27965 14875 27999
rect 15853 27965 15887 27999
rect 16037 27965 16071 27999
rect 17417 27965 17451 27999
rect 18705 27965 18739 27999
rect 23305 27965 23339 27999
rect 24409 27965 24443 27999
rect 25145 27965 25179 27999
rect 27997 27965 28031 27999
rect 28273 27965 28307 27999
rect 34897 27965 34931 27999
rect 11713 27897 11747 27931
rect 31033 27897 31067 27931
rect 1593 27829 1627 27863
rect 13645 27829 13679 27863
rect 20453 27829 20487 27863
rect 22109 27829 22143 27863
rect 23857 27829 23891 27863
rect 25789 27829 25823 27863
rect 26525 27829 26559 27863
rect 29193 27829 29227 27863
rect 32505 27829 32539 27863
rect 36645 27829 36679 27863
rect 16116 27625 16150 27659
rect 28917 27625 28951 27659
rect 35633 27625 35667 27659
rect 7297 27557 7331 27591
rect 18889 27557 18923 27591
rect 23489 27557 23523 27591
rect 31585 27557 31619 27591
rect 36185 27557 36219 27591
rect 37105 27557 37139 27591
rect 8401 27489 8435 27523
rect 10241 27489 10275 27523
rect 12265 27489 12299 27523
rect 13277 27489 13311 27523
rect 15853 27489 15887 27523
rect 18245 27489 18279 27523
rect 18429 27489 18463 27523
rect 19901 27489 19935 27523
rect 20085 27489 20119 27523
rect 22845 27489 22879 27523
rect 24961 27489 24995 27523
rect 30481 27489 30515 27523
rect 32505 27489 32539 27523
rect 33425 27489 33459 27523
rect 33885 27489 33919 27523
rect 34989 27489 35023 27523
rect 7389 27421 7423 27455
rect 9597 27421 9631 27455
rect 14565 27421 14599 27455
rect 15209 27421 15243 27455
rect 19809 27421 19843 27455
rect 20821 27421 20855 27455
rect 21281 27421 21315 27455
rect 22569 27421 22603 27455
rect 23581 27421 23615 27455
rect 27169 27421 27203 27455
rect 30389 27421 30423 27455
rect 31217 27421 31251 27455
rect 31401 27421 31435 27455
rect 32413 27421 32447 27455
rect 33517 27421 33551 27455
rect 35265 27421 35299 27455
rect 36277 27421 36311 27455
rect 36921 27421 36955 27455
rect 8217 27353 8251 27387
rect 10517 27353 10551 27387
rect 13185 27353 13219 27387
rect 15301 27353 15335 27387
rect 25237 27353 25271 27387
rect 27445 27353 27479 27387
rect 7849 27285 7883 27319
rect 8309 27285 8343 27319
rect 9781 27285 9815 27319
rect 12725 27285 12759 27319
rect 13093 27285 13127 27319
rect 14381 27285 14415 27319
rect 17601 27285 17635 27319
rect 18521 27285 18555 27319
rect 19441 27285 19475 27319
rect 20637 27285 20671 27319
rect 21373 27285 21407 27319
rect 22201 27285 22235 27319
rect 22661 27285 22695 27319
rect 26709 27285 26743 27319
rect 30757 27285 30791 27319
rect 32781 27285 32815 27319
rect 35173 27285 35207 27319
rect 9137 27081 9171 27115
rect 9597 27081 9631 27115
rect 11713 27081 11747 27115
rect 12173 27081 12207 27115
rect 15485 27081 15519 27115
rect 24685 27081 24719 27115
rect 25145 27081 25179 27115
rect 25605 27081 25639 27115
rect 26433 27081 26467 27115
rect 28733 27081 28767 27115
rect 30757 27081 30791 27115
rect 10057 27013 10091 27047
rect 12081 27013 12115 27047
rect 13553 27013 13587 27047
rect 19441 27013 19475 27047
rect 22845 27013 22879 27047
rect 23673 27013 23707 27047
rect 24777 27013 24811 27047
rect 33425 27013 33459 27047
rect 9965 26945 9999 26979
rect 11161 26945 11195 26979
rect 15853 26945 15887 26979
rect 17049 26945 17083 26979
rect 20269 26945 20303 26979
rect 22201 26945 22235 26979
rect 25789 26945 25823 26979
rect 26249 26945 26283 26979
rect 27169 26945 27203 26979
rect 28365 26945 28399 26979
rect 28549 26945 28583 26979
rect 29193 26945 29227 26979
rect 30665 26945 30699 26979
rect 31585 26945 31619 26979
rect 32505 26945 32539 26979
rect 33333 26945 33367 26979
rect 34621 26945 34655 26979
rect 35817 26945 35851 26979
rect 36461 26945 36495 26979
rect 36645 26945 36679 26979
rect 7389 26877 7423 26911
rect 7665 26877 7699 26911
rect 10241 26877 10275 26911
rect 12357 26877 12391 26911
rect 13277 26877 13311 26911
rect 15025 26877 15059 26911
rect 15945 26877 15979 26911
rect 16129 26877 16163 26911
rect 19717 26877 19751 26911
rect 21005 26877 21039 26911
rect 24593 26877 24627 26911
rect 27353 26877 27387 26911
rect 30573 26877 30607 26911
rect 32413 26877 32447 26911
rect 34437 26877 34471 26911
rect 34529 26877 34563 26911
rect 35725 26877 35759 26911
rect 31125 26809 31159 26843
rect 36553 26809 36587 26843
rect 11069 26741 11103 26775
rect 17141 26741 17175 26775
rect 17969 26741 18003 26775
rect 22017 26741 22051 26775
rect 29285 26741 29319 26775
rect 31769 26741 31803 26775
rect 32781 26741 32815 26775
rect 34989 26741 35023 26775
rect 35541 26741 35575 26775
rect 7757 26537 7791 26571
rect 8493 26537 8527 26571
rect 16313 26537 16347 26571
rect 18889 26537 18923 26571
rect 22477 26537 22511 26571
rect 27169 26537 27203 26571
rect 28733 26537 28767 26571
rect 30205 26537 30239 26571
rect 34253 26537 34287 26571
rect 37059 26537 37093 26571
rect 11345 26469 11379 26503
rect 16773 26469 16807 26503
rect 23949 26469 23983 26503
rect 26617 26469 26651 26503
rect 10333 26401 10367 26435
rect 11805 26401 11839 26435
rect 12081 26401 12115 26435
rect 13553 26401 13587 26435
rect 14933 26401 14967 26435
rect 15117 26401 15151 26435
rect 17417 26401 17451 26435
rect 18245 26401 18279 26435
rect 18429 26401 18463 26435
rect 19993 26401 20027 26435
rect 20085 26401 20119 26435
rect 20729 26401 20763 26435
rect 23397 26401 23431 26435
rect 26065 26401 26099 26435
rect 31677 26401 31711 26435
rect 32689 26401 32723 26435
rect 33885 26401 33919 26435
rect 35265 26401 35299 26435
rect 35633 26401 35667 26435
rect 7941 26333 7975 26367
rect 8401 26333 8435 26367
rect 10057 26333 10091 26367
rect 11161 26333 11195 26367
rect 16129 26333 16163 26367
rect 17141 26333 17175 26367
rect 17233 26333 17267 26367
rect 23581 26333 23615 26367
rect 24777 26333 24811 26367
rect 25421 26333 25455 26367
rect 27261 26333 27295 26367
rect 27905 26333 27939 26367
rect 31953 26333 31987 26367
rect 32965 26333 32999 26367
rect 33149 26333 33183 26367
rect 33977 26333 34011 26367
rect 14841 26265 14875 26299
rect 21005 26265 21039 26299
rect 25329 26265 25363 26299
rect 28549 26265 28583 26299
rect 28749 26265 28783 26299
rect 32827 26265 32861 26299
rect 33057 26265 33091 26299
rect 9689 26197 9723 26231
rect 10149 26197 10183 26231
rect 14473 26197 14507 26231
rect 18521 26197 18555 26231
rect 19533 26197 19567 26231
rect 19901 26197 19935 26231
rect 23489 26197 23523 26231
rect 24593 26197 24627 26231
rect 26157 26197 26191 26231
rect 26249 26197 26283 26231
rect 27721 26197 27755 26231
rect 28917 26197 28951 26231
rect 33333 26197 33367 26231
rect 15669 25993 15703 26027
rect 19257 25993 19291 26027
rect 26065 25993 26099 26027
rect 26157 25993 26191 26027
rect 30481 25993 30515 26027
rect 33517 25993 33551 26027
rect 14197 25925 14231 25959
rect 18337 25925 18371 25959
rect 19993 25925 20027 25959
rect 27445 25925 27479 25959
rect 30573 25925 30607 25959
rect 33425 25925 33459 25959
rect 8401 25857 8435 25891
rect 9229 25857 9263 25891
rect 12173 25857 12207 25891
rect 13277 25857 13311 25891
rect 16129 25857 16163 25891
rect 19073 25857 19107 25891
rect 22109 25857 22143 25891
rect 24869 25857 24903 25891
rect 24961 25857 24995 25891
rect 29561 25857 29595 25891
rect 29653 25857 29687 25891
rect 29837 25857 29871 25891
rect 30389 25857 30423 25891
rect 30665 25857 30699 25891
rect 31125 25857 31159 25891
rect 31309 25857 31343 25891
rect 32505 25857 32539 25891
rect 32597 25857 32631 25891
rect 32781 25857 32815 25891
rect 33333 25857 33367 25891
rect 33793 25857 33827 25891
rect 9505 25789 9539 25823
rect 13921 25789 13955 25823
rect 18613 25789 18647 25823
rect 19717 25789 19751 25823
rect 22385 25789 22419 25823
rect 25145 25789 25179 25823
rect 26249 25789 26283 25823
rect 27169 25789 27203 25823
rect 36185 25789 36219 25823
rect 36461 25789 36495 25823
rect 10977 25721 11011 25755
rect 23857 25721 23891 25755
rect 29745 25721 29779 25755
rect 32321 25721 32355 25755
rect 34713 25721 34747 25755
rect 8493 25653 8527 25687
rect 12265 25653 12299 25687
rect 13461 25653 13495 25687
rect 16313 25653 16347 25687
rect 16865 25653 16899 25687
rect 21465 25653 21499 25687
rect 24501 25653 24535 25687
rect 25697 25653 25731 25687
rect 28917 25653 28951 25687
rect 29377 25653 29411 25687
rect 31217 25653 31251 25687
rect 32781 25653 32815 25687
rect 8585 25449 8619 25483
rect 12909 25449 12943 25483
rect 18337 25449 18371 25483
rect 19441 25449 19475 25483
rect 20913 25449 20947 25483
rect 28365 25449 28399 25483
rect 31493 25449 31527 25483
rect 31769 25449 31803 25483
rect 32597 25449 32631 25483
rect 35909 25449 35943 25483
rect 36461 25449 36495 25483
rect 9873 25313 9907 25347
rect 11161 25313 11195 25347
rect 14565 25313 14599 25347
rect 16865 25313 16899 25347
rect 19901 25313 19935 25347
rect 20085 25313 20119 25347
rect 23765 25313 23799 25347
rect 23857 25313 23891 25347
rect 24685 25313 24719 25347
rect 26617 25313 26651 25347
rect 30573 25313 30607 25347
rect 31493 25313 31527 25347
rect 33609 25313 33643 25347
rect 7941 25245 7975 25279
rect 8401 25245 8435 25279
rect 10517 25245 10551 25279
rect 14289 25245 14323 25279
rect 16589 25245 16623 25279
rect 21005 25245 21039 25279
rect 22661 25245 22695 25279
rect 23673 25245 23707 25279
rect 24961 25245 24995 25279
rect 25789 25245 25823 25279
rect 29745 25245 29779 25279
rect 30389 25245 30423 25279
rect 30481 25245 30515 25279
rect 31401 25245 31435 25279
rect 32229 25245 32263 25279
rect 34069 25245 34103 25279
rect 34253 25245 34287 25279
rect 35081 25245 35115 25279
rect 35173 25245 35207 25279
rect 35725 25245 35759 25279
rect 36369 25245 36403 25279
rect 11437 25177 11471 25211
rect 26893 25177 26927 25211
rect 32413 25177 32447 25211
rect 33241 25177 33275 25211
rect 33425 25177 33459 25211
rect 34161 25177 34195 25211
rect 7757 25109 7791 25143
rect 9321 25109 9355 25143
rect 9689 25109 9723 25143
rect 9781 25109 9815 25143
rect 10701 25109 10735 25143
rect 16037 25109 16071 25143
rect 19809 25109 19843 25143
rect 22477 25109 22511 25143
rect 23305 25109 23339 25143
rect 24869 25109 24903 25143
rect 25329 25109 25363 25143
rect 25881 25109 25915 25143
rect 34897 25109 34931 25143
rect 10701 24905 10735 24939
rect 12081 24905 12115 24939
rect 21097 24905 21131 24939
rect 23765 24905 23799 24939
rect 25973 24905 26007 24939
rect 27169 24905 27203 24939
rect 29009 24905 29043 24939
rect 30113 24905 30147 24939
rect 34805 24905 34839 24939
rect 7757 24837 7791 24871
rect 10793 24837 10827 24871
rect 13277 24837 13311 24871
rect 19073 24837 19107 24871
rect 21005 24837 21039 24871
rect 22293 24837 22327 24871
rect 29101 24837 29135 24871
rect 9781 24769 9815 24803
rect 9873 24769 9907 24803
rect 14933 24769 14967 24803
rect 15485 24769 15519 24803
rect 15577 24769 15611 24803
rect 16129 24769 16163 24803
rect 17325 24769 17359 24803
rect 17969 24769 18003 24803
rect 19165 24769 19199 24803
rect 20177 24769 20211 24803
rect 26617 24769 26651 24803
rect 27353 24769 27387 24803
rect 27813 24769 27847 24803
rect 27905 24769 27939 24803
rect 28917 24769 28951 24803
rect 29745 24769 29779 24803
rect 30573 24769 30607 24803
rect 31309 24769 31343 24803
rect 31401 24769 31435 24803
rect 32781 24769 32815 24803
rect 32965 24769 32999 24803
rect 33793 24769 33827 24803
rect 36369 24769 36403 24803
rect 36461 24769 36495 24803
rect 7481 24701 7515 24735
rect 10517 24701 10551 24735
rect 12173 24701 12207 24735
rect 12357 24701 12391 24735
rect 13001 24701 13035 24735
rect 13185 24701 13219 24735
rect 14841 24701 14875 24735
rect 17049 24701 17083 24735
rect 19257 24701 19291 24735
rect 21281 24701 21315 24735
rect 22017 24701 22051 24735
rect 24225 24701 24259 24735
rect 24501 24701 24535 24735
rect 29837 24701 29871 24735
rect 33609 24701 33643 24735
rect 34529 24701 34563 24735
rect 34713 24701 34747 24735
rect 11713 24633 11747 24667
rect 17877 24633 17911 24667
rect 20637 24633 20671 24667
rect 26433 24633 26467 24667
rect 28733 24633 28767 24667
rect 29285 24633 29319 24667
rect 9229 24565 9263 24599
rect 11161 24565 11195 24599
rect 13645 24565 13679 24599
rect 16313 24565 16347 24599
rect 18705 24565 18739 24599
rect 19993 24565 20027 24599
rect 29929 24565 29963 24599
rect 30665 24565 30699 24599
rect 33149 24565 33183 24599
rect 33977 24565 34011 24599
rect 35173 24565 35207 24599
rect 7849 24361 7883 24395
rect 15669 24361 15703 24395
rect 20361 24361 20395 24395
rect 23673 24361 23707 24395
rect 27077 24361 27111 24395
rect 32781 24293 32815 24327
rect 8309 24225 8343 24259
rect 8493 24225 8527 24259
rect 10057 24225 10091 24259
rect 12725 24225 12759 24259
rect 17141 24225 17175 24259
rect 17417 24225 17451 24259
rect 19717 24225 19751 24259
rect 19901 24225 19935 24259
rect 25697 24225 25731 24259
rect 26433 24225 26467 24259
rect 31493 24225 31527 24259
rect 31769 24225 31803 24259
rect 32321 24225 32355 24259
rect 33793 24225 33827 24259
rect 34161 24225 34195 24259
rect 35449 24225 35483 24259
rect 1777 24157 1811 24191
rect 7389 24157 7423 24191
rect 11345 24157 11379 24191
rect 13553 24157 13587 24191
rect 14473 24157 14507 24191
rect 15025 24157 15059 24191
rect 18337 24157 18371 24191
rect 21281 24157 21315 24191
rect 23121 24157 23155 24191
rect 23765 24157 23799 24191
rect 25513 24157 25547 24191
rect 26617 24157 26651 24191
rect 26709 24157 26743 24191
rect 29009 24157 29043 24191
rect 29101 24157 29135 24191
rect 32413 24157 32447 24191
rect 33701 24157 33735 24191
rect 36921 24157 36955 24191
rect 8217 24089 8251 24123
rect 10885 24089 10919 24123
rect 11989 24089 12023 24123
rect 29745 24089 29779 24123
rect 35357 24089 35391 24123
rect 1593 24021 1627 24055
rect 7297 24021 7331 24055
rect 11529 24021 11563 24055
rect 13369 24021 13403 24055
rect 14381 24021 14415 24055
rect 15209 24021 15243 24055
rect 18153 24021 18187 24055
rect 19993 24021 20027 24055
rect 21189 24021 21223 24055
rect 22937 24021 22971 24055
rect 25145 24021 25179 24055
rect 25605 24021 25639 24055
rect 33517 24021 33551 24055
rect 34897 24021 34931 24055
rect 35265 24021 35299 24055
rect 37105 24021 37139 24055
rect 9597 23817 9631 23851
rect 10793 23817 10827 23851
rect 10885 23817 10919 23851
rect 12173 23817 12207 23851
rect 14749 23817 14783 23851
rect 16957 23817 16991 23851
rect 19257 23817 19291 23851
rect 24041 23817 24075 23851
rect 24409 23817 24443 23851
rect 26157 23817 26191 23851
rect 28917 23817 28951 23851
rect 32873 23817 32907 23851
rect 36829 23817 36863 23851
rect 12081 23749 12115 23783
rect 13277 23749 13311 23783
rect 17785 23749 17819 23783
rect 19993 23749 20027 23783
rect 13001 23681 13035 23715
rect 15393 23681 15427 23715
rect 17049 23681 17083 23715
rect 22845 23681 22879 23715
rect 24501 23681 24535 23715
rect 29745 23681 29779 23715
rect 32505 23681 32539 23715
rect 33517 23681 33551 23715
rect 34437 23681 34471 23715
rect 35081 23681 35115 23715
rect 7021 23613 7055 23647
rect 7297 23613 7331 23647
rect 8769 23613 8803 23647
rect 9689 23613 9723 23647
rect 9781 23613 9815 23647
rect 10977 23613 11011 23647
rect 11989 23613 12023 23647
rect 15669 23613 15703 23647
rect 17509 23613 17543 23647
rect 19717 23613 19751 23647
rect 23121 23613 23155 23647
rect 24685 23613 24719 23647
rect 25881 23613 25915 23647
rect 26065 23613 26099 23647
rect 27169 23613 27203 23647
rect 27445 23613 27479 23647
rect 30113 23613 30147 23647
rect 32413 23613 32447 23647
rect 33609 23613 33643 23647
rect 33885 23613 33919 23647
rect 35357 23613 35391 23647
rect 34621 23545 34655 23579
rect 9229 23477 9263 23511
rect 10425 23477 10459 23511
rect 12541 23477 12575 23511
rect 21465 23477 21499 23511
rect 26525 23477 26559 23511
rect 31539 23477 31573 23511
rect 6193 23273 6227 23307
rect 9137 23273 9171 23307
rect 12725 23273 12759 23307
rect 14381 23273 14415 23307
rect 18613 23273 18647 23307
rect 19533 23273 19567 23307
rect 26525 23273 26559 23307
rect 27813 23273 27847 23307
rect 29009 23273 29043 23307
rect 30481 23273 30515 23307
rect 31677 23273 31711 23307
rect 33425 23273 33459 23307
rect 33609 23273 33643 23307
rect 35173 23273 35207 23307
rect 12265 23205 12299 23239
rect 6837 23137 6871 23171
rect 8401 23137 8435 23171
rect 9689 23137 9723 23171
rect 10517 23137 10551 23171
rect 13185 23137 13219 23171
rect 13277 23137 13311 23171
rect 15853 23137 15887 23171
rect 16129 23137 16163 23171
rect 19993 23137 20027 23171
rect 20177 23137 20211 23171
rect 21649 23137 21683 23171
rect 22293 23137 22327 23171
rect 24041 23137 24075 23171
rect 25605 23137 25639 23171
rect 36921 23137 36955 23171
rect 6009 23069 6043 23103
rect 8309 23069 8343 23103
rect 9505 23069 9539 23103
rect 13093 23069 13127 23103
rect 16773 23069 16807 23103
rect 17233 23069 17267 23103
rect 18521 23069 18555 23103
rect 21465 23069 21499 23103
rect 25421 23069 25455 23103
rect 26341 23069 26375 23103
rect 27721 23069 27755 23103
rect 28733 23069 28767 23103
rect 28825 23069 28859 23103
rect 29745 23069 29779 23103
rect 29929 23069 29963 23103
rect 30389 23069 30423 23103
rect 33609 23069 33643 23103
rect 33793 23069 33827 23103
rect 7021 23001 7055 23035
rect 10793 23001 10827 23035
rect 21373 23001 21407 23035
rect 22569 23001 22603 23035
rect 28457 23001 28491 23035
rect 32965 23001 32999 23035
rect 36645 23001 36679 23035
rect 6929 22933 6963 22967
rect 7389 22933 7423 22967
rect 7849 22933 7883 22967
rect 8217 22933 8251 22967
rect 9597 22933 9631 22967
rect 16681 22933 16715 22967
rect 17325 22933 17359 22967
rect 19901 22933 19935 22967
rect 21005 22933 21039 22967
rect 25053 22933 25087 22967
rect 25513 22933 25547 22967
rect 28641 22933 28675 22967
rect 29837 22933 29871 22967
rect 8401 22729 8435 22763
rect 10885 22729 10919 22763
rect 13461 22729 13495 22763
rect 25329 22729 25363 22763
rect 26341 22729 26375 22763
rect 28917 22729 28951 22763
rect 35909 22729 35943 22763
rect 36461 22729 36495 22763
rect 11989 22661 12023 22695
rect 14933 22661 14967 22695
rect 27445 22661 27479 22695
rect 30665 22661 30699 22695
rect 32689 22661 32723 22695
rect 32807 22661 32841 22695
rect 33517 22661 33551 22695
rect 35265 22661 35299 22695
rect 6653 22593 6687 22627
rect 9137 22593 9171 22627
rect 11713 22593 11747 22627
rect 13921 22593 13955 22627
rect 16129 22593 16163 22627
rect 18613 22593 18647 22627
rect 19349 22593 19383 22627
rect 20545 22593 20579 22627
rect 22017 22593 22051 22627
rect 22753 22593 22787 22627
rect 26157 22593 26191 22627
rect 29929 22593 29963 22627
rect 30573 22593 30607 22627
rect 30757 22593 30791 22627
rect 32505 22593 32539 22627
rect 32597 22593 32631 22627
rect 35725 22593 35759 22627
rect 36553 22593 36587 22627
rect 6929 22525 6963 22559
rect 9413 22525 9447 22559
rect 18337 22525 18371 22559
rect 20637 22525 20671 22559
rect 20729 22525 20763 22559
rect 23029 22525 23063 22559
rect 24501 22525 24535 22559
rect 25421 22525 25455 22559
rect 25513 22525 25547 22559
rect 27169 22525 27203 22559
rect 30113 22525 30147 22559
rect 32965 22525 32999 22559
rect 15209 22457 15243 22491
rect 16313 22457 16347 22491
rect 14105 22389 14139 22423
rect 16865 22389 16899 22423
rect 19257 22389 19291 22423
rect 20177 22389 20211 22423
rect 22109 22389 22143 22423
rect 24961 22389 24995 22423
rect 29745 22389 29779 22423
rect 32321 22389 32355 22423
rect 7297 22185 7331 22219
rect 9505 22185 9539 22219
rect 10793 22185 10827 22219
rect 14546 22185 14580 22219
rect 31953 22185 31987 22219
rect 8033 22049 8067 22083
rect 10057 22049 10091 22083
rect 11989 22049 12023 22083
rect 13093 22049 13127 22083
rect 17601 22049 17635 22083
rect 18337 22049 18371 22083
rect 20361 22049 20395 22083
rect 23305 22049 23339 22083
rect 25697 22049 25731 22083
rect 27629 22049 27663 22083
rect 28733 22049 28767 22083
rect 30021 22049 30055 22083
rect 30297 22049 30331 22083
rect 31401 22049 31435 22083
rect 32321 22049 32355 22083
rect 35265 22049 35299 22083
rect 36829 22049 36863 22083
rect 7481 21981 7515 22015
rect 8125 21981 8159 22015
rect 9321 21981 9355 22015
rect 9965 21981 9999 22015
rect 10609 21981 10643 22015
rect 12081 21981 12115 22015
rect 12909 21981 12943 22015
rect 14289 21981 14323 22015
rect 16773 21981 16807 22015
rect 18429 21981 18463 22015
rect 19717 21981 19751 22015
rect 23213 21981 23247 22015
rect 24041 21981 24075 22015
rect 24777 21981 24811 22015
rect 25973 21981 26007 22015
rect 27077 21981 27111 22015
rect 27537 21981 27571 22015
rect 28825 21981 28859 22015
rect 29929 21981 29963 22015
rect 31125 21981 31159 22015
rect 31217 21981 31251 22015
rect 32229 21981 32263 22015
rect 33609 21981 33643 22015
rect 33793 21981 33827 22015
rect 33977 21981 34011 22015
rect 35081 21981 35115 22015
rect 36001 21981 36035 22015
rect 36737 21981 36771 22015
rect 17325 21913 17359 21947
rect 20637 21913 20671 21947
rect 25881 21913 25915 21947
rect 33701 21913 33735 21947
rect 12541 21845 12575 21879
rect 13001 21845 13035 21879
rect 16037 21845 16071 21879
rect 16681 21845 16715 21879
rect 18521 21845 18555 21879
rect 18889 21845 18923 21879
rect 19901 21845 19935 21879
rect 22109 21845 22143 21879
rect 23857 21845 23891 21879
rect 24685 21845 24719 21879
rect 26341 21845 26375 21879
rect 26985 21845 27019 21879
rect 29193 21845 29227 21879
rect 33425 21845 33459 21879
rect 34897 21845 34931 21879
rect 36093 21845 36127 21879
rect 12081 21641 12115 21675
rect 13921 21641 13955 21675
rect 14749 21641 14783 21675
rect 18245 21641 18279 21675
rect 20453 21641 20487 21675
rect 20913 21641 20947 21675
rect 22477 21641 22511 21675
rect 23673 21641 23707 21675
rect 25605 21641 25639 21675
rect 25697 21641 25731 21675
rect 28917 21641 28951 21675
rect 29561 21641 29595 21675
rect 30481 21641 30515 21675
rect 32873 21641 32907 21675
rect 13553 21573 13587 21607
rect 29377 21573 29411 21607
rect 7849 21505 7883 21539
rect 10149 21505 10183 21539
rect 12173 21505 12207 21539
rect 14657 21505 14691 21539
rect 15853 21505 15887 21539
rect 17325 21505 17359 21539
rect 19993 21505 20027 21539
rect 20821 21505 20855 21539
rect 22385 21505 22419 21539
rect 23581 21505 23615 21539
rect 24409 21505 24443 21539
rect 26433 21505 26467 21539
rect 27169 21505 27203 21539
rect 29653 21505 29687 21539
rect 32505 21505 32539 21539
rect 33793 21505 33827 21539
rect 13277 21437 13311 21471
rect 13461 21437 13495 21471
rect 16129 21437 16163 21471
rect 17601 21437 17635 21471
rect 19717 21437 19751 21471
rect 21005 21437 21039 21471
rect 22569 21437 22603 21471
rect 25789 21437 25823 21471
rect 27445 21437 27479 21471
rect 30297 21437 30331 21471
rect 30389 21437 30423 21471
rect 32413 21437 32447 21471
rect 33701 21437 33735 21471
rect 34989 21437 35023 21471
rect 35265 21437 35299 21471
rect 22017 21369 22051 21403
rect 26617 21369 26651 21403
rect 29377 21369 29411 21403
rect 7941 21301 7975 21335
rect 9965 21301 9999 21335
rect 24317 21301 24351 21335
rect 25237 21301 25271 21335
rect 30849 21301 30883 21335
rect 34069 21301 34103 21335
rect 36737 21301 36771 21335
rect 8585 21097 8619 21131
rect 26525 21097 26559 21131
rect 28733 21097 28767 21131
rect 32965 21097 32999 21131
rect 6837 20961 6871 20995
rect 9689 20961 9723 20995
rect 12633 20961 12667 20995
rect 19625 20961 19659 20995
rect 22385 20961 22419 20995
rect 23305 20961 23339 20995
rect 25145 20961 25179 20995
rect 25881 20961 25915 20995
rect 29101 20961 29135 20995
rect 30205 20961 30239 20995
rect 33517 20961 33551 20995
rect 35357 20961 35391 20995
rect 35449 20961 35483 20995
rect 9505 20893 9539 20927
rect 10977 20893 11011 20927
rect 11437 20893 11471 20927
rect 12449 20893 12483 20927
rect 14289 20893 14323 20927
rect 15393 20893 15427 20927
rect 17693 20893 17727 20927
rect 23029 20893 23063 20927
rect 24961 20893 24995 20927
rect 27261 20893 27295 20927
rect 29009 20893 29043 20927
rect 32689 20893 32723 20927
rect 32781 20893 32815 20927
rect 32965 20893 32999 20927
rect 35265 20893 35299 20927
rect 7113 20825 7147 20859
rect 17417 20825 17451 20859
rect 18521 20825 18555 20859
rect 21373 20825 21407 20859
rect 22201 20825 22235 20859
rect 27537 20825 27571 20859
rect 30481 20825 30515 20859
rect 33701 20825 33735 20859
rect 9137 20757 9171 20791
rect 9597 20757 9631 20791
rect 10885 20757 10919 20791
rect 11621 20757 11655 20791
rect 12081 20757 12115 20791
rect 12541 20757 12575 20791
rect 14473 20757 14507 20791
rect 15301 20757 15335 20791
rect 15945 20757 15979 20791
rect 18797 20757 18831 20791
rect 21833 20757 21867 20791
rect 22293 20757 22327 20791
rect 24593 20757 24627 20791
rect 25053 20757 25087 20791
rect 26065 20757 26099 20791
rect 26157 20757 26191 20791
rect 31953 20757 31987 20791
rect 33793 20757 33827 20791
rect 34161 20757 34195 20791
rect 34897 20757 34931 20791
rect 7389 20553 7423 20587
rect 8401 20553 8435 20587
rect 11161 20553 11195 20587
rect 13461 20553 13495 20587
rect 15853 20553 15887 20587
rect 17049 20553 17083 20587
rect 19717 20553 19751 20587
rect 24777 20553 24811 20587
rect 25605 20553 25639 20587
rect 25697 20553 25731 20587
rect 27537 20553 27571 20587
rect 29837 20553 29871 20587
rect 30205 20553 30239 20587
rect 30665 20553 30699 20587
rect 32413 20553 32447 20587
rect 35173 20553 35207 20587
rect 9689 20485 9723 20519
rect 11989 20485 12023 20519
rect 14381 20485 14415 20519
rect 1777 20417 1811 20451
rect 7573 20417 7607 20451
rect 8493 20417 8527 20451
rect 9413 20417 9447 20451
rect 11713 20417 11747 20451
rect 16865 20417 16899 20451
rect 17693 20417 17727 20451
rect 18613 20417 18647 20451
rect 19625 20417 19659 20451
rect 20637 20417 20671 20451
rect 21281 20417 21315 20451
rect 22569 20417 22603 20451
rect 26433 20417 26467 20451
rect 28549 20417 28583 20451
rect 30849 20417 30883 20451
rect 31493 20417 31527 20451
rect 32505 20417 32539 20451
rect 33517 20417 33551 20451
rect 34529 20417 34563 20451
rect 34989 20417 35023 20451
rect 35817 20417 35851 20451
rect 36737 20417 36771 20451
rect 8677 20349 8711 20383
rect 14105 20349 14139 20383
rect 19809 20349 19843 20383
rect 23029 20349 23063 20383
rect 23305 20349 23339 20383
rect 25789 20349 25823 20383
rect 27629 20349 27663 20383
rect 27721 20349 27755 20383
rect 29653 20349 29687 20383
rect 29745 20349 29779 20383
rect 33425 20349 33459 20383
rect 33885 20349 33919 20383
rect 1593 20281 1627 20315
rect 8033 20281 8067 20315
rect 19257 20281 19291 20315
rect 27169 20281 27203 20315
rect 36921 20281 36955 20315
rect 17601 20213 17635 20247
rect 18797 20213 18831 20247
rect 20821 20213 20855 20247
rect 21373 20213 21407 20247
rect 22385 20213 22419 20247
rect 25237 20213 25271 20247
rect 26617 20213 26651 20247
rect 28457 20213 28491 20247
rect 31309 20213 31343 20247
rect 34345 20213 34379 20247
rect 35725 20213 35759 20247
rect 9873 20009 9907 20043
rect 12449 20009 12483 20043
rect 14289 20009 14323 20043
rect 19625 20009 19659 20043
rect 22201 20009 22235 20043
rect 23305 20009 23339 20043
rect 24593 20009 24627 20043
rect 28457 20009 28491 20043
rect 32597 20009 32631 20043
rect 10517 19873 10551 19907
rect 11529 19873 11563 19907
rect 11713 19873 11747 19907
rect 13093 19873 13127 19907
rect 13277 19873 13311 19907
rect 14841 19873 14875 19907
rect 16313 19873 16347 19907
rect 20453 19873 20487 19907
rect 23949 19873 23983 19907
rect 25605 19873 25639 19907
rect 26985 19873 27019 19907
rect 31585 19873 31619 19907
rect 34069 19873 34103 19907
rect 34345 19873 34379 19907
rect 8585 19805 8619 19839
rect 9321 19805 9355 19839
rect 10241 19805 10275 19839
rect 12357 19805 12391 19839
rect 13369 19805 13403 19839
rect 14657 19805 14691 19839
rect 15669 19805 15703 19839
rect 18705 19805 18739 19839
rect 19441 19805 19475 19839
rect 23673 19805 23707 19839
rect 24777 19805 24811 19839
rect 26709 19805 26743 19839
rect 10333 19737 10367 19771
rect 11437 19737 11471 19771
rect 14749 19737 14783 19771
rect 16589 19737 16623 19771
rect 20729 19737 20763 19771
rect 31309 19737 31343 19771
rect 8401 19669 8435 19703
rect 9229 19669 9263 19703
rect 11069 19669 11103 19703
rect 13737 19669 13771 19703
rect 15853 19669 15887 19703
rect 18061 19669 18095 19703
rect 18797 19669 18831 19703
rect 23765 19669 23799 19703
rect 25789 19669 25823 19703
rect 25881 19669 25915 19703
rect 26249 19669 26283 19703
rect 29837 19669 29871 19703
rect 10241 19465 10275 19499
rect 10609 19465 10643 19499
rect 13001 19465 13035 19499
rect 13369 19465 13403 19499
rect 16865 19465 16899 19499
rect 17233 19465 17267 19499
rect 20637 19465 20671 19499
rect 21005 19465 21039 19499
rect 23857 19465 23891 19499
rect 24961 19465 24995 19499
rect 25789 19465 25823 19499
rect 26157 19465 26191 19499
rect 28917 19465 28951 19499
rect 30849 19465 30883 19499
rect 21097 19397 21131 19431
rect 22385 19397 22419 19431
rect 25053 19397 25087 19431
rect 29469 19397 29503 19431
rect 8033 19329 8067 19363
rect 10701 19329 10735 19363
rect 11897 19329 11931 19363
rect 12357 19329 12391 19363
rect 13461 19329 13495 19363
rect 14565 19329 14599 19363
rect 19901 19329 19935 19363
rect 22109 19329 22143 19363
rect 27169 19329 27203 19363
rect 29561 19329 29595 19363
rect 30941 19329 30975 19363
rect 34069 19329 34103 19363
rect 8309 19261 8343 19295
rect 9781 19261 9815 19295
rect 10793 19261 10827 19295
rect 13553 19261 13587 19295
rect 14841 19261 14875 19295
rect 17325 19261 17359 19295
rect 17417 19261 17451 19295
rect 19625 19261 19659 19295
rect 21189 19261 21223 19295
rect 25145 19261 25179 19295
rect 26249 19261 26283 19295
rect 26341 19261 26375 19295
rect 27445 19261 27479 19295
rect 33793 19261 33827 19295
rect 16313 19193 16347 19227
rect 11713 19125 11747 19159
rect 12541 19125 12575 19159
rect 18153 19125 18187 19159
rect 24593 19125 24627 19159
rect 32321 19125 32355 19159
rect 7757 18921 7791 18955
rect 12081 18921 12115 18955
rect 13737 18921 13771 18955
rect 14381 18921 14415 18955
rect 17049 18921 17083 18955
rect 18797 18921 18831 18955
rect 19441 18921 19475 18955
rect 26341 18921 26375 18955
rect 26985 18921 27019 18955
rect 31033 18921 31067 18955
rect 32873 18921 32907 18955
rect 6009 18785 6043 18819
rect 9137 18785 9171 18819
rect 11437 18785 11471 18819
rect 11621 18785 11655 18819
rect 15577 18785 15611 18819
rect 17693 18785 17727 18819
rect 21189 18785 21223 18819
rect 24593 18785 24627 18819
rect 30757 18785 30791 18819
rect 32137 18785 32171 18819
rect 12909 18717 12943 18751
rect 13553 18717 13587 18751
rect 14289 18717 14323 18751
rect 15301 18717 15335 18751
rect 15393 18717 15427 18751
rect 16497 18717 16531 18751
rect 17417 18717 17451 18751
rect 18889 18717 18923 18751
rect 22109 18717 22143 18751
rect 22845 18717 22879 18751
rect 23857 18717 23891 18751
rect 26801 18717 26835 18751
rect 27629 18717 27663 18751
rect 29009 18717 29043 18751
rect 29193 18717 29227 18751
rect 29837 18717 29871 18751
rect 30021 18717 30055 18751
rect 30665 18717 30699 18751
rect 32321 18717 32355 18751
rect 32781 18717 32815 18751
rect 35081 18717 35115 18751
rect 6285 18649 6319 18683
rect 9413 18649 9447 18683
rect 20913 18649 20947 18683
rect 21833 18649 21867 18683
rect 24869 18649 24903 18683
rect 28365 18649 28399 18683
rect 10885 18581 10919 18615
rect 11713 18581 11747 18615
rect 13001 18581 13035 18615
rect 14933 18581 14967 18615
rect 16221 18581 16255 18615
rect 17509 18581 17543 18615
rect 22937 18581 22971 18615
rect 24041 18581 24075 18615
rect 29009 18581 29043 18615
rect 29929 18581 29963 18615
rect 34989 18581 35023 18615
rect 6009 18377 6043 18411
rect 7205 18377 7239 18411
rect 8217 18377 8251 18411
rect 11161 18377 11195 18411
rect 14841 18377 14875 18411
rect 15209 18377 15243 18411
rect 19073 18377 19107 18411
rect 19441 18377 19475 18411
rect 20821 18377 20855 18411
rect 24317 18377 24351 18411
rect 31769 18377 31803 18411
rect 32505 18377 32539 18411
rect 12909 18309 12943 18343
rect 17141 18309 17175 18343
rect 25237 18309 25271 18343
rect 27445 18309 27479 18343
rect 28825 18309 28859 18343
rect 30297 18309 30331 18343
rect 32321 18309 32355 18343
rect 33149 18309 33183 18343
rect 5825 18241 5859 18275
rect 7297 18241 7331 18275
rect 8125 18241 8159 18275
rect 8769 18241 8803 18275
rect 9413 18241 9447 18275
rect 11989 18241 12023 18275
rect 16129 18241 16163 18275
rect 19533 18241 19567 18275
rect 20729 18241 20763 18275
rect 24225 18241 24259 18275
rect 26065 18241 26099 18275
rect 27169 18241 27203 18275
rect 28549 18241 28583 18275
rect 28642 18241 28676 18275
rect 28917 18241 28951 18275
rect 29055 18241 29089 18275
rect 30021 18241 30055 18275
rect 32597 18241 32631 18275
rect 33241 18241 33275 18275
rect 33793 18241 33827 18275
rect 9689 18173 9723 18207
rect 12633 18173 12667 18207
rect 14381 18173 14415 18207
rect 15301 18173 15335 18207
rect 15485 18173 15519 18207
rect 16865 18173 16899 18207
rect 19717 18173 19751 18207
rect 21005 18173 21039 18207
rect 22017 18173 22051 18207
rect 22293 18173 22327 18207
rect 25329 18173 25363 18207
rect 25513 18173 25547 18207
rect 34069 18173 34103 18207
rect 8953 18105 8987 18139
rect 16313 18105 16347 18139
rect 32321 18105 32355 18139
rect 12081 18037 12115 18071
rect 18613 18037 18647 18071
rect 20361 18037 20395 18071
rect 23765 18037 23799 18071
rect 24869 18037 24903 18071
rect 26249 18037 26283 18071
rect 29193 18037 29227 18071
rect 35541 18037 35575 18071
rect 8217 17833 8251 17867
rect 9597 17833 9631 17867
rect 13093 17833 13127 17867
rect 22569 17833 22603 17867
rect 25973 17833 26007 17867
rect 28641 17833 28675 17867
rect 33977 17833 34011 17867
rect 6469 17765 6503 17799
rect 16037 17765 16071 17799
rect 20729 17765 20763 17799
rect 35173 17765 35207 17799
rect 7113 17697 7147 17731
rect 10701 17697 10735 17731
rect 11345 17697 11379 17731
rect 14841 17697 14875 17731
rect 15025 17697 15059 17731
rect 16957 17697 16991 17731
rect 17141 17697 17175 17731
rect 18245 17697 18279 17731
rect 18429 17697 18463 17731
rect 20085 17697 20119 17731
rect 23673 17697 23707 17731
rect 23857 17697 23891 17731
rect 25329 17697 25363 17731
rect 25513 17697 25547 17731
rect 26709 17697 26743 17731
rect 30021 17697 30055 17731
rect 31217 17697 31251 17731
rect 33517 17697 33551 17731
rect 5825 17629 5859 17663
rect 8033 17629 8067 17663
rect 9505 17629 9539 17663
rect 10609 17629 10643 17663
rect 15117 17629 15151 17663
rect 20361 17629 20395 17663
rect 21373 17629 21407 17663
rect 21925 17629 21959 17663
rect 22753 17629 22787 17663
rect 24593 17629 24627 17663
rect 26433 17629 26467 17663
rect 28825 17629 28859 17663
rect 29009 17629 29043 17663
rect 29929 17629 29963 17663
rect 32965 17629 32999 17663
rect 33609 17629 33643 17663
rect 34897 17629 34931 17663
rect 35633 17629 35667 17663
rect 35817 17629 35851 17663
rect 6837 17561 6871 17595
rect 11621 17561 11655 17595
rect 16313 17561 16347 17595
rect 18521 17561 18555 17595
rect 20269 17561 20303 17595
rect 23581 17561 23615 17595
rect 25605 17561 25639 17595
rect 34989 17561 35023 17595
rect 35173 17561 35207 17595
rect 6009 17493 6043 17527
rect 6929 17493 6963 17527
rect 10149 17493 10183 17527
rect 10517 17493 10551 17527
rect 15485 17493 15519 17527
rect 17233 17493 17267 17527
rect 17601 17493 17635 17527
rect 18889 17493 18923 17527
rect 21189 17493 21223 17527
rect 22017 17493 22051 17527
rect 23213 17493 23247 17527
rect 24777 17493 24811 17527
rect 28181 17493 28215 17527
rect 30297 17493 30331 17527
rect 35725 17493 35759 17527
rect 8309 17289 8343 17323
rect 8769 17289 8803 17323
rect 9137 17289 9171 17323
rect 10425 17289 10459 17323
rect 11713 17289 11747 17323
rect 12173 17289 12207 17323
rect 17233 17289 17267 17323
rect 18889 17289 18923 17323
rect 19717 17289 19751 17323
rect 24593 17289 24627 17323
rect 25421 17289 25455 17323
rect 28273 17289 28307 17323
rect 29469 17289 29503 17323
rect 36645 17289 36679 17323
rect 5917 17221 5951 17255
rect 10333 17221 10367 17255
rect 17325 17221 17359 17255
rect 21189 17221 21223 17255
rect 28825 17221 28859 17255
rect 28917 17221 28951 17255
rect 30297 17221 30331 17255
rect 35173 17221 35207 17255
rect 1777 17153 1811 17187
rect 5825 17153 5859 17187
rect 12081 17153 12115 17187
rect 13185 17153 13219 17187
rect 13277 17153 13311 17187
rect 24685 17153 24719 17187
rect 25789 17153 25823 17187
rect 27353 17153 27387 17187
rect 28549 17153 28583 17187
rect 29561 17153 29595 17187
rect 30021 17153 30055 17187
rect 32321 17153 32355 17187
rect 34897 17153 34931 17187
rect 6561 17085 6595 17119
rect 6837 17085 6871 17119
rect 9229 17085 9263 17119
rect 9321 17085 9355 17119
rect 10609 17085 10643 17119
rect 12357 17085 12391 17119
rect 13093 17085 13127 17119
rect 14565 17085 14599 17119
rect 14841 17085 14875 17119
rect 16313 17085 16347 17119
rect 17417 17085 17451 17119
rect 18613 17085 18647 17119
rect 18797 17085 18831 17119
rect 21465 17085 21499 17119
rect 22017 17085 22051 17119
rect 22293 17085 22327 17119
rect 24869 17085 24903 17119
rect 25881 17085 25915 17119
rect 25973 17085 26007 17119
rect 28457 17085 28491 17119
rect 32597 17085 32631 17119
rect 34069 17085 34103 17119
rect 23765 17017 23799 17051
rect 1593 16949 1627 16983
rect 9965 16949 9999 16983
rect 13645 16949 13679 16983
rect 16865 16949 16899 16983
rect 19257 16949 19291 16983
rect 24225 16949 24259 16983
rect 27261 16949 27295 16983
rect 31769 16949 31803 16983
rect 14381 16745 14415 16779
rect 18613 16745 18647 16779
rect 21189 16745 21223 16779
rect 22293 16745 22327 16779
rect 25770 16745 25804 16779
rect 27261 16745 27295 16779
rect 29837 16745 29871 16779
rect 30757 16745 30791 16779
rect 30941 16745 30975 16779
rect 35081 16745 35115 16779
rect 35265 16745 35299 16779
rect 36001 16745 36035 16779
rect 24961 16677 24995 16711
rect 32597 16677 32631 16711
rect 6837 16609 6871 16643
rect 6929 16609 6963 16643
rect 8033 16609 8067 16643
rect 8217 16609 8251 16643
rect 9137 16609 9171 16643
rect 12725 16609 12759 16643
rect 12909 16609 12943 16643
rect 16865 16609 16899 16643
rect 19441 16609 19475 16643
rect 23489 16609 23523 16643
rect 23581 16609 23615 16643
rect 25513 16609 25547 16643
rect 6745 16541 6779 16575
rect 11621 16541 11655 16575
rect 13645 16541 13679 16575
rect 14657 16541 14691 16575
rect 15485 16541 15519 16575
rect 16129 16541 16163 16575
rect 22109 16541 22143 16575
rect 23397 16541 23431 16575
rect 27813 16541 27847 16575
rect 27905 16541 27939 16575
rect 28457 16541 28491 16575
rect 29745 16541 29779 16575
rect 30021 16541 30055 16575
rect 31677 16541 31711 16575
rect 31769 16541 31803 16575
rect 32689 16541 32723 16575
rect 33149 16541 33183 16575
rect 33241 16541 33275 16575
rect 33977 16541 34011 16575
rect 35909 16541 35943 16575
rect 36921 16541 36955 16575
rect 9413 16473 9447 16507
rect 12633 16473 12667 16507
rect 17141 16473 17175 16507
rect 19717 16473 19751 16507
rect 24685 16473 24719 16507
rect 31125 16473 31159 16507
rect 34897 16473 34931 16507
rect 35113 16473 35147 16507
rect 6377 16405 6411 16439
rect 7573 16405 7607 16439
rect 7941 16405 7975 16439
rect 10885 16405 10919 16439
rect 11713 16405 11747 16439
rect 12265 16405 12299 16439
rect 13461 16405 13495 16439
rect 15669 16405 15703 16439
rect 16221 16405 16255 16439
rect 23029 16405 23063 16439
rect 28549 16405 28583 16439
rect 30297 16405 30331 16439
rect 30915 16405 30949 16439
rect 33885 16405 33919 16439
rect 37105 16405 37139 16439
rect 6929 16201 6963 16235
rect 8125 16201 8159 16235
rect 10241 16201 10275 16235
rect 11713 16201 11747 16235
rect 12081 16201 12115 16235
rect 15669 16201 15703 16235
rect 17141 16201 17175 16235
rect 18061 16201 18095 16235
rect 19073 16201 19107 16235
rect 19717 16201 19751 16235
rect 20361 16201 20395 16235
rect 23397 16201 23431 16235
rect 24225 16201 24259 16235
rect 24593 16201 24627 16235
rect 30021 16201 30055 16235
rect 8953 16133 8987 16167
rect 13553 16133 13587 16167
rect 23489 16133 23523 16167
rect 25697 16133 25731 16167
rect 28641 16133 28675 16167
rect 28733 16133 28767 16167
rect 31401 16133 31435 16167
rect 32597 16133 32631 16167
rect 7021 16065 7055 16099
rect 7941 16065 7975 16099
rect 9045 16065 9079 16099
rect 10149 16065 10183 16099
rect 10977 16065 11011 16099
rect 12173 16065 12207 16099
rect 15577 16065 15611 16099
rect 16957 16065 16991 16099
rect 18153 16065 18187 16099
rect 18889 16065 18923 16099
rect 19625 16065 19659 16099
rect 20269 16065 20303 16099
rect 22385 16065 22419 16099
rect 24685 16065 24719 16099
rect 25789 16065 25823 16099
rect 27353 16065 27387 16099
rect 28365 16065 28399 16099
rect 28458 16065 28492 16099
rect 28871 16065 28905 16099
rect 29469 16065 29503 16099
rect 29561 16065 29595 16099
rect 29745 16065 29779 16099
rect 29837 16065 29871 16099
rect 30665 16065 30699 16099
rect 30849 16065 30883 16099
rect 31309 16065 31343 16099
rect 31493 16065 31527 16099
rect 32413 16065 32447 16099
rect 32689 16065 32723 16099
rect 34069 16065 34103 16099
rect 34713 16065 34747 16099
rect 35357 16065 35391 16099
rect 35541 16065 35575 16099
rect 36185 16065 36219 16099
rect 36645 16065 36679 16099
rect 7205 15997 7239 16031
rect 9137 15997 9171 16031
rect 12265 15997 12299 16031
rect 13277 15997 13311 16031
rect 15025 15997 15059 16031
rect 23581 15997 23615 16031
rect 24777 15997 24811 16031
rect 25513 15997 25547 16031
rect 34529 15997 34563 16031
rect 8585 15929 8619 15963
rect 23029 15929 23063 15963
rect 26157 15929 26191 15963
rect 33977 15929 34011 15963
rect 35357 15929 35391 15963
rect 6561 15861 6595 15895
rect 11161 15861 11195 15895
rect 22201 15861 22235 15895
rect 27261 15861 27295 15895
rect 29009 15861 29043 15895
rect 30849 15861 30883 15895
rect 32413 15861 32447 15895
rect 34897 15861 34931 15895
rect 36093 15861 36127 15895
rect 36737 15861 36771 15895
rect 8033 15657 8067 15691
rect 11510 15657 11544 15691
rect 13001 15657 13035 15691
rect 15209 15657 15243 15691
rect 23397 15657 23431 15691
rect 25053 15657 25087 15691
rect 27905 15657 27939 15691
rect 29193 15657 29227 15691
rect 32597 15657 32631 15691
rect 14473 15589 14507 15623
rect 6285 15521 6319 15555
rect 9689 15521 9723 15555
rect 11253 15521 11287 15555
rect 21925 15521 21959 15555
rect 28733 15521 28767 15555
rect 28825 15521 28859 15555
rect 30389 15521 30423 15555
rect 30665 15521 30699 15555
rect 34345 15521 34379 15555
rect 35357 15521 35391 15555
rect 35633 15521 35667 15555
rect 5825 15453 5859 15487
rect 9505 15453 9539 15487
rect 10517 15453 10551 15487
rect 14657 15453 14691 15487
rect 15393 15453 15427 15487
rect 16313 15453 16347 15487
rect 21649 15453 21683 15487
rect 24777 15453 24811 15487
rect 27353 15453 27387 15487
rect 27813 15453 27847 15487
rect 28457 15453 28491 15487
rect 28641 15453 28675 15487
rect 29009 15453 29043 15487
rect 29745 15453 29779 15487
rect 29929 15453 29963 15487
rect 6561 15385 6595 15419
rect 16037 15385 16071 15419
rect 27077 15385 27111 15419
rect 34069 15385 34103 15419
rect 5733 15317 5767 15351
rect 9137 15317 9171 15351
rect 9597 15317 9631 15351
rect 10425 15317 10459 15351
rect 25605 15317 25639 15351
rect 29837 15317 29871 15351
rect 32137 15317 32171 15351
rect 37105 15317 37139 15351
rect 6009 15113 6043 15147
rect 6653 15113 6687 15147
rect 7113 15113 7147 15147
rect 15301 15113 15335 15147
rect 22661 15113 22695 15147
rect 28365 15113 28399 15147
rect 29193 15113 29227 15147
rect 31125 15113 31159 15147
rect 32489 15113 32523 15147
rect 33241 15113 33275 15147
rect 13369 15045 13403 15079
rect 13737 15045 13771 15079
rect 14473 15045 14507 15079
rect 23213 15045 23247 15079
rect 25697 15045 25731 15079
rect 26525 15045 26559 15079
rect 31677 15045 31711 15079
rect 32689 15045 32723 15079
rect 5825 14977 5859 15011
rect 7021 14977 7055 15011
rect 8309 14977 8343 15011
rect 8953 14977 8987 15011
rect 11713 14977 11747 15011
rect 12725 14977 12759 15011
rect 14749 14977 14783 15011
rect 15393 14977 15427 15011
rect 22569 14977 22603 15011
rect 24593 14977 24627 15011
rect 27537 14977 27571 15011
rect 28549 14977 28583 15011
rect 29331 14977 29365 15011
rect 29469 14977 29503 15011
rect 29561 14977 29595 15011
rect 29689 14977 29723 15011
rect 29837 14977 29871 15011
rect 30941 14977 30975 15011
rect 31769 14977 31803 15011
rect 33333 14977 33367 15011
rect 33885 14977 33919 15011
rect 36277 14977 36311 15011
rect 7205 14909 7239 14943
rect 9229 14909 9263 14943
rect 10701 14909 10735 14943
rect 23949 14909 23983 14943
rect 27629 14909 27663 14943
rect 27721 14909 27755 14943
rect 30757 14909 30791 14943
rect 34161 14909 34195 14943
rect 8493 14841 8527 14875
rect 32321 14841 32355 14875
rect 11897 14773 11931 14807
rect 12449 14773 12483 14807
rect 24777 14773 24811 14807
rect 27169 14773 27203 14807
rect 32505 14773 32539 14807
rect 35633 14773 35667 14807
rect 36185 14773 36219 14807
rect 7849 14569 7883 14603
rect 11713 14569 11747 14603
rect 21189 14569 21223 14603
rect 27721 14569 27755 14603
rect 28181 14569 28215 14603
rect 28641 14569 28675 14603
rect 31585 14569 31619 14603
rect 32413 14569 32447 14603
rect 34253 14569 34287 14603
rect 35541 14569 35575 14603
rect 13185 14501 13219 14535
rect 6101 14433 6135 14467
rect 9781 14433 9815 14467
rect 9873 14433 9907 14467
rect 11069 14433 11103 14467
rect 12265 14433 12299 14467
rect 22937 14433 22971 14467
rect 24961 14433 24995 14467
rect 27445 14433 27479 14467
rect 29929 14433 29963 14467
rect 30389 14433 30423 14467
rect 35173 14433 35207 14467
rect 5457 14365 5491 14399
rect 8401 14365 8435 14399
rect 10885 14365 10919 14399
rect 13461 14365 13495 14399
rect 23581 14365 23615 14399
rect 27353 14365 27387 14399
rect 28365 14365 28399 14399
rect 28457 14365 28491 14399
rect 28733 14365 28767 14399
rect 30021 14365 30055 14399
rect 31033 14365 31067 14399
rect 31677 14365 31711 14399
rect 32229 14365 32263 14399
rect 32413 14365 32447 14399
rect 32873 14365 32907 14399
rect 34069 14365 34103 14399
rect 34253 14365 34287 14399
rect 35265 14365 35299 14399
rect 6377 14297 6411 14331
rect 9689 14297 9723 14331
rect 12173 14297 12207 14331
rect 22661 14297 22695 14331
rect 25237 14297 25271 14331
rect 30297 14297 30331 14331
rect 5641 14229 5675 14263
rect 8585 14229 8619 14263
rect 9321 14229 9355 14263
rect 10517 14229 10551 14263
rect 10977 14229 11011 14263
rect 12081 14229 12115 14263
rect 23397 14229 23431 14263
rect 26709 14229 26743 14263
rect 29745 14229 29779 14263
rect 30941 14229 30975 14263
rect 33057 14229 33091 14263
rect 7021 14025 7055 14059
rect 7481 14025 7515 14059
rect 10057 14025 10091 14059
rect 13829 14025 13863 14059
rect 21373 14025 21407 14059
rect 22477 14025 22511 14059
rect 23305 14025 23339 14059
rect 23673 14025 23707 14059
rect 23765 14025 23799 14059
rect 30297 14025 30331 14059
rect 33241 14025 33275 14059
rect 8585 13957 8619 13991
rect 12357 13957 12391 13991
rect 22385 13957 22419 13991
rect 25145 13957 25179 13991
rect 29653 13957 29687 13991
rect 7389 13889 7423 13923
rect 8309 13889 8343 13923
rect 10517 13889 10551 13923
rect 14289 13889 14323 13923
rect 21465 13889 21499 13923
rect 24869 13889 24903 13923
rect 27261 13889 27295 13923
rect 28733 13889 28767 13923
rect 28825 13889 28859 13923
rect 29009 13889 29043 13923
rect 29101 13889 29135 13923
rect 29561 13889 29595 13923
rect 30205 13889 30239 13923
rect 31033 13889 31067 13923
rect 31493 13889 31527 13923
rect 32873 13889 32907 13923
rect 33793 13889 33827 13923
rect 7665 13821 7699 13855
rect 12081 13821 12115 13855
rect 14381 13821 14415 13855
rect 22293 13821 22327 13855
rect 23949 13821 23983 13855
rect 26617 13821 26651 13855
rect 27537 13821 27571 13855
rect 32597 13821 32631 13855
rect 32781 13821 32815 13855
rect 22845 13753 22879 13787
rect 28549 13753 28583 13787
rect 10701 13685 10735 13719
rect 30849 13685 30883 13719
rect 31677 13685 31711 13719
rect 33885 13685 33919 13719
rect 7297 13481 7331 13515
rect 9137 13481 9171 13515
rect 12081 13481 12115 13515
rect 24593 13481 24627 13515
rect 26157 13481 26191 13515
rect 27077 13481 27111 13515
rect 31493 13481 31527 13515
rect 33701 13481 33735 13515
rect 8493 13413 8527 13447
rect 22477 13413 22511 13447
rect 24041 13413 24075 13447
rect 9781 13345 9815 13379
rect 10333 13345 10367 13379
rect 10609 13345 10643 13379
rect 23121 13345 23155 13379
rect 25145 13345 25179 13379
rect 28825 13345 28859 13379
rect 29745 13345 29779 13379
rect 1777 13277 1811 13311
rect 6561 13277 6595 13311
rect 7389 13277 7423 13311
rect 8585 13277 8619 13311
rect 9505 13277 9539 13311
rect 9597 13277 9631 13311
rect 13461 13277 13495 13311
rect 14381 13277 14415 13311
rect 21925 13277 21959 13311
rect 23857 13277 23891 13311
rect 31953 13277 31987 13311
rect 34345 13277 34379 13311
rect 36921 13277 36955 13311
rect 12725 13209 12759 13243
rect 25881 13209 25915 13243
rect 28549 13209 28583 13243
rect 30021 13209 30055 13243
rect 32229 13209 32263 13243
rect 34253 13209 34287 13243
rect 1593 13141 1627 13175
rect 6653 13141 6687 13175
rect 14473 13141 14507 13175
rect 21741 13141 21775 13175
rect 22845 13141 22879 13175
rect 22937 13141 22971 13175
rect 24961 13141 24995 13175
rect 25053 13141 25087 13175
rect 37105 13141 37139 13175
rect 9505 12937 9539 12971
rect 10425 12937 10459 12971
rect 10793 12937 10827 12971
rect 10885 12937 10919 12971
rect 14289 12937 14323 12971
rect 23213 12937 23247 12971
rect 23673 12937 23707 12971
rect 25881 12937 25915 12971
rect 27261 12937 27295 12971
rect 28273 12937 28307 12971
rect 28825 12937 28859 12971
rect 30573 12937 30607 12971
rect 31769 12937 31803 12971
rect 34529 12937 34563 12971
rect 12081 12869 12115 12903
rect 24777 12869 24811 12903
rect 31309 12869 31343 12903
rect 33057 12869 33091 12903
rect 6561 12801 6595 12835
rect 13461 12801 13495 12835
rect 13737 12801 13771 12835
rect 14381 12801 14415 12835
rect 17785 12801 17819 12835
rect 22109 12801 22143 12835
rect 23581 12801 23615 12835
rect 25973 12801 26007 12835
rect 27353 12801 27387 12835
rect 28181 12801 28215 12835
rect 29009 12801 29043 12835
rect 30205 12801 30239 12835
rect 31401 12801 31435 12835
rect 32781 12801 32815 12835
rect 6837 12733 6871 12767
rect 9597 12733 9631 12767
rect 9781 12733 9815 12767
rect 10977 12733 11011 12767
rect 12173 12733 12207 12767
rect 12357 12733 12391 12767
rect 17601 12733 17635 12767
rect 23857 12733 23891 12767
rect 24869 12733 24903 12767
rect 25053 12733 25087 12767
rect 29929 12733 29963 12767
rect 30113 12733 30147 12767
rect 31217 12733 31251 12767
rect 8309 12597 8343 12631
rect 9137 12597 9171 12631
rect 11713 12597 11747 12631
rect 22201 12597 22235 12631
rect 24409 12597 24443 12631
rect 6377 12393 6411 12427
rect 8585 12393 8619 12427
rect 13553 12393 13587 12427
rect 22845 12393 22879 12427
rect 26709 12393 26743 12427
rect 31585 12393 31619 12427
rect 6837 12257 6871 12291
rect 9689 12257 9723 12291
rect 11805 12257 11839 12291
rect 21097 12257 21131 12291
rect 23949 12257 23983 12291
rect 24961 12257 24995 12291
rect 27169 12257 27203 12291
rect 32045 12257 32079 12291
rect 32137 12257 32171 12291
rect 33333 12257 33367 12291
rect 6193 12189 6227 12223
rect 9505 12189 9539 12223
rect 10517 12189 10551 12223
rect 11161 12189 11195 12223
rect 14473 12189 14507 12223
rect 23673 12189 23707 12223
rect 28917 12189 28951 12223
rect 29929 12189 29963 12223
rect 30573 12189 30607 12223
rect 34161 12189 34195 12223
rect 34897 12189 34931 12223
rect 7113 12121 7147 12155
rect 12081 12121 12115 12155
rect 14381 12121 14415 12155
rect 21373 12121 21407 12155
rect 25237 12121 25271 12155
rect 28641 12121 28675 12155
rect 30481 12121 30515 12155
rect 33149 12121 33183 12155
rect 9137 12053 9171 12087
rect 9597 12053 9631 12087
rect 10609 12053 10643 12087
rect 11345 12053 11379 12087
rect 23305 12053 23339 12087
rect 23765 12053 23799 12087
rect 29745 12053 29779 12087
rect 31953 12053 31987 12087
rect 32781 12053 32815 12087
rect 33241 12053 33275 12087
rect 33977 12053 34011 12087
rect 34989 12053 35023 12087
rect 6561 11849 6595 11883
rect 7849 11849 7883 11883
rect 9413 11849 9447 11883
rect 9505 11849 9539 11883
rect 10701 11849 10735 11883
rect 24593 11849 24627 11883
rect 28457 11849 28491 11883
rect 29101 11849 29135 11883
rect 30021 11849 30055 11883
rect 31401 11849 31435 11883
rect 34805 11849 34839 11883
rect 13737 11781 13771 11815
rect 27537 11781 27571 11815
rect 31309 11781 31343 11815
rect 6929 11713 6963 11747
rect 7757 11713 7791 11747
rect 8401 11713 8435 11747
rect 10793 11713 10827 11747
rect 12633 11713 12667 11747
rect 13461 11713 13495 11747
rect 22017 11713 22051 11747
rect 25789 11713 25823 11747
rect 27445 11713 27479 11747
rect 28549 11713 28583 11747
rect 29193 11713 29227 11747
rect 30113 11713 30147 11747
rect 32505 11713 32539 11747
rect 7021 11645 7055 11679
rect 7205 11645 7239 11679
rect 9689 11645 9723 11679
rect 10609 11645 10643 11679
rect 11805 11645 11839 11679
rect 22293 11645 22327 11679
rect 23765 11645 23799 11679
rect 24685 11645 24719 11679
rect 24777 11645 24811 11679
rect 25881 11645 25915 11679
rect 25973 11645 26007 11679
rect 27353 11645 27387 11679
rect 29929 11645 29963 11679
rect 31217 11645 31251 11679
rect 33057 11645 33091 11679
rect 33333 11645 33367 11679
rect 9045 11577 9079 11611
rect 27905 11577 27939 11611
rect 30481 11577 30515 11611
rect 8585 11509 8619 11543
rect 11161 11509 11195 11543
rect 24225 11509 24259 11543
rect 25421 11509 25455 11543
rect 31769 11509 31803 11543
rect 32413 11509 32447 11543
rect 7665 11305 7699 11339
rect 11897 11305 11931 11339
rect 12357 11305 12391 11339
rect 22293 11305 22327 11339
rect 23029 11305 23063 11339
rect 24041 11305 24075 11339
rect 25329 11305 25363 11339
rect 29837 11305 29871 11339
rect 31327 11305 31361 11339
rect 33793 11237 33827 11271
rect 12817 11169 12851 11203
rect 12909 11169 12943 11203
rect 24777 11169 24811 11203
rect 24869 11169 24903 11203
rect 26893 11169 26927 11203
rect 27629 11169 27663 11203
rect 31585 11169 31619 11203
rect 32045 11169 32079 11203
rect 6561 11101 6595 11135
rect 7849 11101 7883 11135
rect 9505 11101 9539 11135
rect 10149 11101 10183 11135
rect 13737 11101 13771 11135
rect 22477 11101 22511 11135
rect 22937 11101 22971 11135
rect 23857 11101 23891 11135
rect 35081 11101 35115 11135
rect 10425 11033 10459 11067
rect 13645 11033 13679 11067
rect 24961 11033 24995 11067
rect 26617 11033 26651 11067
rect 26709 11033 26743 11067
rect 27721 11033 27755 11067
rect 27813 11033 27847 11067
rect 28733 11033 28767 11067
rect 29101 11033 29135 11067
rect 32321 11033 32355 11067
rect 34989 11033 35023 11067
rect 6377 10965 6411 10999
rect 9597 10965 9631 10999
rect 12725 10965 12759 10999
rect 26249 10965 26283 10999
rect 28181 10965 28215 10999
rect 10241 10761 10275 10795
rect 10701 10761 10735 10795
rect 24685 10761 24719 10795
rect 25881 10761 25915 10795
rect 30297 10761 30331 10795
rect 30757 10761 30791 10795
rect 32505 10761 32539 10795
rect 33425 10761 33459 10795
rect 34253 10761 34287 10795
rect 8769 10693 8803 10727
rect 27445 10693 27479 10727
rect 29561 10693 29595 10727
rect 6929 10625 6963 10659
rect 7941 10625 7975 10659
rect 8493 10625 8527 10659
rect 10885 10625 10919 10659
rect 12173 10625 12207 10659
rect 17877 10625 17911 10659
rect 22753 10625 22787 10659
rect 23581 10625 23615 10659
rect 24961 10625 24995 10659
rect 27169 10625 27203 10659
rect 29837 10625 29871 10659
rect 30665 10625 30699 10659
rect 31677 10625 31711 10659
rect 32321 10625 32355 10659
rect 33333 10625 33367 10659
rect 34345 10625 34379 10659
rect 7021 10557 7055 10591
rect 7205 10557 7239 10591
rect 12449 10557 12483 10591
rect 17693 10557 17727 10591
rect 25973 10557 26007 10591
rect 26157 10557 26191 10591
rect 28089 10557 28123 10591
rect 30849 10557 30883 10591
rect 33517 10557 33551 10591
rect 6561 10489 6595 10523
rect 32965 10489 32999 10523
rect 7849 10421 7883 10455
rect 13921 10421 13955 10455
rect 22569 10421 22603 10455
rect 23305 10421 23339 10455
rect 25513 10421 25547 10455
rect 31493 10421 31527 10455
rect 11805 10217 11839 10251
rect 24041 10217 24075 10251
rect 28917 10217 28951 10251
rect 29745 10217 29779 10251
rect 31309 10217 31343 10251
rect 33333 10217 33367 10251
rect 26341 10149 26375 10183
rect 6101 10081 6135 10115
rect 9137 10081 9171 10115
rect 12725 10081 12759 10115
rect 12909 10081 12943 10115
rect 22293 10081 22327 10115
rect 24593 10081 24627 10115
rect 28365 10081 28399 10115
rect 30297 10081 30331 10115
rect 32689 10081 32723 10115
rect 8401 10013 8435 10047
rect 11621 10013 11655 10047
rect 12633 10013 12667 10047
rect 27537 10013 27571 10047
rect 29101 10013 29135 10047
rect 30113 10013 30147 10047
rect 33517 10013 33551 10047
rect 34161 10013 34195 10047
rect 6377 9945 6411 9979
rect 9413 9945 9447 9979
rect 22569 9945 22603 9979
rect 24869 9945 24903 9979
rect 31033 9945 31067 9979
rect 32505 9945 32539 9979
rect 7849 9877 7883 9911
rect 8585 9877 8619 9911
rect 10885 9877 10919 9911
rect 12265 9877 12299 9911
rect 30205 9877 30239 9911
rect 32137 9877 32171 9911
rect 32597 9877 32631 9911
rect 33977 9877 34011 9911
rect 8493 9673 8527 9707
rect 10057 9673 10091 9707
rect 13461 9673 13495 9707
rect 14381 9673 14415 9707
rect 28733 9673 28767 9707
rect 28825 9673 28859 9707
rect 8861 9605 8895 9639
rect 10149 9605 10183 9639
rect 23765 9605 23799 9639
rect 25513 9605 25547 9639
rect 27629 9605 27663 9639
rect 30297 9605 30331 9639
rect 33149 9605 33183 9639
rect 1777 9537 1811 9571
rect 7389 9537 7423 9571
rect 7481 9537 7515 9571
rect 10977 9537 11011 9571
rect 11713 9537 11747 9571
rect 14289 9537 14323 9571
rect 22661 9537 22695 9571
rect 23857 9537 23891 9571
rect 24961 9537 24995 9571
rect 25421 9537 25455 9571
rect 26065 9537 26099 9571
rect 27537 9537 27571 9571
rect 30021 9537 30055 9571
rect 36737 9537 36771 9571
rect 7665 9469 7699 9503
rect 8953 9469 8987 9503
rect 9045 9469 9079 9503
rect 10241 9469 10275 9503
rect 11989 9469 12023 9503
rect 14565 9469 14599 9503
rect 22845 9469 22879 9503
rect 27721 9469 27755 9503
rect 28917 9469 28951 9503
rect 32873 9469 32907 9503
rect 7021 9401 7055 9435
rect 11161 9401 11195 9435
rect 24777 9401 24811 9435
rect 28365 9401 28399 9435
rect 1593 9333 1627 9367
rect 9689 9333 9723 9367
rect 13921 9333 13955 9367
rect 26157 9333 26191 9367
rect 27169 9333 27203 9367
rect 31769 9333 31803 9367
rect 34621 9333 34655 9367
rect 36921 9333 36955 9367
rect 10793 9129 10827 9163
rect 12081 9129 12115 9163
rect 26433 9129 26467 9163
rect 31401 9129 31435 9163
rect 33333 9129 33367 9163
rect 33977 9129 34011 9163
rect 10241 9061 10275 9095
rect 6837 8993 6871 9027
rect 8401 8993 8435 9027
rect 9689 8993 9723 9027
rect 12725 8993 12759 9027
rect 24685 8993 24719 9027
rect 26893 8993 26927 9027
rect 30573 8993 30607 9027
rect 32045 8993 32079 9027
rect 32689 8993 32723 9027
rect 6193 8925 6227 8959
rect 8217 8925 8251 8959
rect 9873 8925 9907 8959
rect 10885 8925 10919 8959
rect 11529 8925 11563 8959
rect 12449 8925 12483 8959
rect 13553 8925 13587 8959
rect 14289 8925 14323 8959
rect 29745 8925 29779 8959
rect 31769 8925 31803 8959
rect 32965 8925 32999 8959
rect 33885 8925 33919 8959
rect 7021 8857 7055 8891
rect 9781 8857 9815 8891
rect 12541 8857 12575 8891
rect 14565 8857 14599 8891
rect 24961 8857 24995 8891
rect 27169 8857 27203 8891
rect 31861 8857 31895 8891
rect 32873 8857 32907 8891
rect 6101 8789 6135 8823
rect 6929 8789 6963 8823
rect 7389 8789 7423 8823
rect 7849 8789 7883 8823
rect 8309 8789 8343 8823
rect 11345 8789 11379 8823
rect 13645 8789 13679 8823
rect 16037 8789 16071 8823
rect 28641 8789 28675 8823
rect 9413 8585 9447 8619
rect 12081 8585 12115 8619
rect 13645 8585 13679 8619
rect 15853 8585 15887 8619
rect 26525 8585 26559 8619
rect 27813 8585 27847 8619
rect 30481 8585 30515 8619
rect 31677 8585 31711 8619
rect 32689 8585 32723 8619
rect 33517 8585 33551 8619
rect 33885 8585 33919 8619
rect 33977 8585 34011 8619
rect 10885 8517 10919 8551
rect 15761 8517 15795 8551
rect 25053 8517 25087 8551
rect 5825 8449 5859 8483
rect 11989 8449 12023 8483
rect 13461 8449 13495 8483
rect 14473 8449 14507 8483
rect 14565 8449 14599 8483
rect 25789 8449 25823 8483
rect 26433 8449 26467 8483
rect 27905 8449 27939 8483
rect 28733 8449 28767 8483
rect 31125 8449 31159 8483
rect 31769 8449 31803 8483
rect 34897 8449 34931 8483
rect 8033 8381 8067 8415
rect 8309 8381 8343 8415
rect 11161 8381 11195 8415
rect 14657 8381 14691 8415
rect 15577 8381 15611 8415
rect 16865 8381 16899 8415
rect 17141 8381 17175 8415
rect 27721 8381 27755 8415
rect 29009 8381 29043 8415
rect 32505 8381 32539 8415
rect 32597 8381 32631 8415
rect 34069 8381 34103 8415
rect 6009 8313 6043 8347
rect 6561 8313 6595 8347
rect 14105 8313 14139 8347
rect 18613 8313 18647 8347
rect 30941 8313 30975 8347
rect 33057 8313 33091 8347
rect 34805 8313 34839 8347
rect 16221 8245 16255 8279
rect 28273 8245 28307 8279
rect 6745 8041 6779 8075
rect 10701 8041 10735 8075
rect 15117 8041 15151 8075
rect 16497 8041 16531 8075
rect 17325 8041 17359 8075
rect 25329 8041 25363 8075
rect 27169 8041 27203 8075
rect 30481 8041 30515 8075
rect 31296 8041 31330 8075
rect 34897 8041 34931 8075
rect 28365 7973 28399 8007
rect 7205 7905 7239 7939
rect 7297 7905 7331 7939
rect 13645 7905 13679 7939
rect 15577 7905 15611 7939
rect 15669 7905 15703 7939
rect 28917 7905 28951 7939
rect 29929 7905 29963 7939
rect 30021 7905 30055 7939
rect 31033 7905 31067 7939
rect 33333 7905 33367 7939
rect 7941 7837 7975 7871
rect 9321 7837 9355 7871
rect 10793 7837 10827 7871
rect 14289 7837 14323 7871
rect 16313 7837 16347 7871
rect 17233 7837 17267 7871
rect 25513 7837 25547 7871
rect 27353 7837 27387 7871
rect 28733 7837 28767 7871
rect 30113 7837 30147 7871
rect 33609 7837 33643 7871
rect 35081 7837 35115 7871
rect 7113 7769 7147 7803
rect 12817 7769 12851 7803
rect 8125 7701 8159 7735
rect 9229 7701 9263 7735
rect 14381 7701 14415 7735
rect 15485 7701 15519 7735
rect 28825 7701 28859 7735
rect 32781 7701 32815 7735
rect 33517 7701 33551 7735
rect 33977 7701 34011 7735
rect 7481 7497 7515 7531
rect 15761 7497 15795 7531
rect 31309 7497 31343 7531
rect 34529 7497 34563 7531
rect 8953 7429 8987 7463
rect 15025 7429 15059 7463
rect 9229 7361 9263 7395
rect 12357 7361 12391 7395
rect 12817 7361 12851 7395
rect 15945 7361 15979 7395
rect 27353 7361 27387 7395
rect 27997 7361 28031 7395
rect 31401 7361 31435 7395
rect 15301 7293 15335 7327
rect 30481 7293 30515 7327
rect 30757 7293 30791 7327
rect 32781 7293 32815 7327
rect 33057 7293 33091 7327
rect 12173 7157 12207 7191
rect 12909 7157 12943 7191
rect 13553 7157 13587 7191
rect 27169 7157 27203 7191
rect 27905 7157 27939 7191
rect 29009 7157 29043 7191
rect 12068 6953 12102 6987
rect 26512 6953 26546 6987
rect 15393 6817 15427 6851
rect 29009 6817 29043 6851
rect 29837 6817 29871 6851
rect 31125 6817 31159 6851
rect 32229 6817 32263 6851
rect 33425 6817 33459 6851
rect 11805 6749 11839 6783
rect 16221 6749 16255 6783
rect 16865 6749 16899 6783
rect 26249 6749 26283 6783
rect 32505 6749 32539 6783
rect 33333 6749 33367 6783
rect 34161 6749 34195 6783
rect 28825 6681 28859 6715
rect 30021 6681 30055 6715
rect 31217 6681 31251 6715
rect 32413 6681 32447 6715
rect 13553 6613 13587 6647
rect 16681 6613 16715 6647
rect 27997 6613 28031 6647
rect 28457 6613 28491 6647
rect 28917 6613 28951 6647
rect 30113 6613 30147 6647
rect 30481 6613 30515 6647
rect 31309 6613 31343 6647
rect 31677 6613 31711 6647
rect 32873 6613 32907 6647
rect 33977 6613 34011 6647
rect 12633 6409 12667 6443
rect 13093 6409 13127 6443
rect 14657 6409 14691 6443
rect 16221 6409 16255 6443
rect 27169 6409 27203 6443
rect 27537 6409 27571 6443
rect 29009 6409 29043 6443
rect 31217 6409 31251 6443
rect 11989 6273 12023 6307
rect 13001 6273 13035 6307
rect 14749 6273 14783 6307
rect 15853 6273 15887 6307
rect 16865 6273 16899 6307
rect 26617 6273 26651 6307
rect 28549 6273 28583 6307
rect 31401 6273 31435 6307
rect 35081 6273 35115 6307
rect 13277 6205 13311 6239
rect 14841 6205 14875 6239
rect 15577 6205 15611 6239
rect 15761 6205 15795 6239
rect 27629 6205 27663 6239
rect 27813 6205 27847 6239
rect 30481 6205 30515 6239
rect 30757 6205 30791 6239
rect 32689 6205 32723 6239
rect 32965 6205 32999 6239
rect 34897 6137 34931 6171
rect 11805 6069 11839 6103
rect 14289 6069 14323 6103
rect 16957 6069 16991 6103
rect 26433 6069 26467 6103
rect 28457 6069 28491 6103
rect 34437 6069 34471 6103
rect 15025 5865 15059 5899
rect 27813 5865 27847 5899
rect 29101 5865 29135 5899
rect 30113 5865 30147 5899
rect 33885 5865 33919 5899
rect 11621 5729 11655 5763
rect 14473 5729 14507 5763
rect 14565 5729 14599 5763
rect 15853 5729 15887 5763
rect 16129 5729 16163 5763
rect 26341 5729 26375 5763
rect 30941 5729 30975 5763
rect 33241 5729 33275 5763
rect 1777 5661 1811 5695
rect 11345 5661 11379 5695
rect 13553 5661 13587 5695
rect 14657 5661 14691 5695
rect 26065 5661 26099 5695
rect 29009 5661 29043 5695
rect 30021 5661 30055 5695
rect 33517 5661 33551 5695
rect 36921 5661 36955 5695
rect 31217 5593 31251 5627
rect 1593 5525 1627 5559
rect 13093 5525 13127 5559
rect 13737 5525 13771 5559
rect 17601 5525 17635 5559
rect 32689 5525 32723 5559
rect 33425 5525 33459 5559
rect 37105 5525 37139 5559
rect 11069 5321 11103 5355
rect 13369 5321 13403 5355
rect 27261 5321 27295 5355
rect 27721 5321 27755 5355
rect 30389 5321 30423 5355
rect 31585 5321 31619 5355
rect 32689 5321 32723 5355
rect 33793 5321 33827 5355
rect 15301 5253 15335 5287
rect 29561 5253 29595 5287
rect 32781 5253 32815 5287
rect 10517 5185 10551 5219
rect 10977 5185 11011 5219
rect 11989 5185 12023 5219
rect 13001 5185 13035 5219
rect 15577 5185 15611 5219
rect 16221 5185 16255 5219
rect 17049 5185 17083 5219
rect 18429 5185 18463 5219
rect 27629 5185 27663 5219
rect 28549 5185 28583 5219
rect 30757 5185 30791 5219
rect 30849 5185 30883 5219
rect 31769 5185 31803 5219
rect 33701 5185 33735 5219
rect 12725 5117 12759 5151
rect 12909 5117 12943 5151
rect 13829 5117 13863 5151
rect 27905 5117 27939 5151
rect 29653 5117 29687 5151
rect 29837 5117 29871 5151
rect 30941 5117 30975 5151
rect 32873 5117 32907 5151
rect 10425 4981 10459 5015
rect 12081 4981 12115 5015
rect 16129 4981 16163 5015
rect 16865 4981 16899 5015
rect 18337 4981 18371 5015
rect 28733 4981 28767 5015
rect 29193 4981 29227 5015
rect 32321 4981 32355 5015
rect 12173 4777 12207 4811
rect 13645 4777 13679 4811
rect 14289 4777 14323 4811
rect 31953 4777 31987 4811
rect 32689 4777 32723 4811
rect 10977 4709 11011 4743
rect 22477 4709 22511 4743
rect 31493 4709 31527 4743
rect 11621 4641 11655 4675
rect 12817 4641 12851 4675
rect 14749 4641 14783 4675
rect 14841 4641 14875 4675
rect 16497 4641 16531 4675
rect 18613 4641 18647 4675
rect 23121 4641 23155 4675
rect 28733 4641 28767 4675
rect 30021 4641 30055 4675
rect 10333 4573 10367 4607
rect 13553 4573 13587 4607
rect 17141 4573 17175 4607
rect 19993 4573 20027 4607
rect 20637 4573 20671 4607
rect 21833 4573 21867 4607
rect 27721 4573 27755 4607
rect 28549 4573 28583 4607
rect 29745 4573 29779 4607
rect 32137 4573 32171 4607
rect 32781 4573 32815 4607
rect 11345 4505 11379 4539
rect 16405 4505 16439 4539
rect 17417 4505 17451 4539
rect 22845 4505 22879 4539
rect 10517 4437 10551 4471
rect 11437 4437 11471 4471
rect 12541 4437 12575 4471
rect 12633 4437 12667 4471
rect 14657 4437 14691 4471
rect 15945 4437 15979 4471
rect 16313 4437 16347 4471
rect 18061 4437 18095 4471
rect 18429 4437 18463 4471
rect 18521 4437 18555 4471
rect 19809 4437 19843 4471
rect 20545 4437 20579 4471
rect 22017 4437 22051 4471
rect 22937 4437 22971 4471
rect 27537 4437 27571 4471
rect 28181 4437 28215 4471
rect 28641 4437 28675 4471
rect 12449 4233 12483 4267
rect 12909 4233 12943 4267
rect 18889 4233 18923 4267
rect 24593 4233 24627 4267
rect 29469 4233 29503 4267
rect 29837 4233 29871 4267
rect 10793 4165 10827 4199
rect 13737 4165 13771 4199
rect 19625 4165 19659 4199
rect 22293 4165 22327 4199
rect 27537 4165 27571 4199
rect 12541 4097 12575 4131
rect 16313 4097 16347 4131
rect 30665 4097 30699 4131
rect 30757 4097 30791 4131
rect 10885 4029 10919 4063
rect 11069 4029 11103 4063
rect 12357 4029 12391 4063
rect 13829 4029 13863 4063
rect 14013 4029 14047 4063
rect 14565 4029 14599 4063
rect 16037 4029 16071 4063
rect 17141 4029 17175 4063
rect 17417 4029 17451 4063
rect 19349 4029 19383 4063
rect 22017 4029 22051 4063
rect 23765 4029 23799 4063
rect 24685 4029 24719 4063
rect 24777 4029 24811 4063
rect 27261 4029 27295 4063
rect 29009 4029 29043 4063
rect 29929 4029 29963 4063
rect 30021 4029 30055 4063
rect 13369 3961 13403 3995
rect 24225 3961 24259 3995
rect 10425 3893 10459 3927
rect 21097 3893 21131 3927
rect 12265 3689 12299 3723
rect 16313 3689 16347 3723
rect 17509 3689 17543 3723
rect 18153 3689 18187 3723
rect 23765 3689 23799 3723
rect 28089 3689 28123 3723
rect 15485 3621 15519 3655
rect 22477 3621 22511 3655
rect 10517 3553 10551 3587
rect 13369 3553 13403 3587
rect 14841 3553 14875 3587
rect 16957 3553 16991 3587
rect 18797 3553 18831 3587
rect 20269 3553 20303 3587
rect 23121 3553 23155 3587
rect 28917 3553 28951 3587
rect 9873 3485 9907 3519
rect 15025 3485 15059 3519
rect 17693 3485 17727 3519
rect 22845 3485 22879 3519
rect 23857 3485 23891 3519
rect 24777 3485 24811 3519
rect 27997 3485 28031 3519
rect 28641 3485 28675 3519
rect 10793 3417 10827 3451
rect 16773 3417 16807 3451
rect 18521 3417 18555 3451
rect 20545 3417 20579 3451
rect 10057 3349 10091 3383
rect 12725 3349 12759 3383
rect 13093 3349 13127 3383
rect 13185 3349 13219 3383
rect 15117 3349 15151 3383
rect 16681 3349 16715 3383
rect 18613 3349 18647 3383
rect 22017 3349 22051 3383
rect 22937 3349 22971 3383
rect 24685 3349 24719 3383
rect 11161 3145 11195 3179
rect 14105 3145 14139 3179
rect 19901 3145 19935 3179
rect 20361 3145 20395 3179
rect 12633 3077 12667 3111
rect 16037 3077 16071 3111
rect 20729 3077 20763 3111
rect 22569 3077 22603 3111
rect 1777 3009 1811 3043
rect 10977 3009 11011 3043
rect 11713 3009 11747 3043
rect 16313 3009 16347 3043
rect 17141 3009 17175 3043
rect 19717 3009 19751 3043
rect 20821 3009 20855 3043
rect 22845 3009 22879 3043
rect 25053 3009 25087 3043
rect 36737 3009 36771 3043
rect 12357 2941 12391 2975
rect 17417 2941 17451 2975
rect 21005 2941 21039 2975
rect 24777 2941 24811 2975
rect 11897 2873 11931 2907
rect 23305 2873 23339 2907
rect 1593 2805 1627 2839
rect 14565 2805 14599 2839
rect 18889 2805 18923 2839
rect 36921 2805 36955 2839
rect 10517 2601 10551 2635
rect 14933 2601 14967 2635
rect 15485 2601 15519 2635
rect 16313 2601 16347 2635
rect 18705 2601 18739 2635
rect 20085 2601 20119 2635
rect 22109 2601 22143 2635
rect 24777 2601 24811 2635
rect 25237 2601 25271 2635
rect 32551 2601 32585 2635
rect 34897 2601 34931 2635
rect 11713 2533 11747 2567
rect 13461 2465 13495 2499
rect 17877 2465 17911 2499
rect 18061 2465 18095 2499
rect 20545 2465 20579 2499
rect 20637 2465 20671 2499
rect 22937 2465 22971 2499
rect 1777 2397 1811 2431
rect 4445 2397 4479 2431
rect 7205 2397 7239 2431
rect 9873 2397 9907 2431
rect 10333 2397 10367 2431
rect 11161 2397 11195 2431
rect 14841 2397 14875 2431
rect 15669 2397 15703 2431
rect 16129 2397 16163 2431
rect 18613 2397 18647 2431
rect 19625 2397 19659 2431
rect 21465 2397 21499 2431
rect 22201 2397 22235 2431
rect 23213 2397 23247 2431
rect 24593 2397 24627 2431
rect 25421 2397 25455 2431
rect 32321 2397 32355 2431
rect 35081 2397 35115 2431
rect 36737 2397 36771 2431
rect 11069 2329 11103 2363
rect 13185 2329 13219 2363
rect 17785 2329 17819 2363
rect 23121 2329 23155 2363
rect 29837 2329 29871 2363
rect 1593 2261 1627 2295
rect 4261 2261 4295 2295
rect 7021 2261 7055 2295
rect 9689 2261 9723 2295
rect 17417 2261 17451 2295
rect 19441 2261 19475 2295
rect 20453 2261 20487 2295
rect 21281 2261 21315 2295
rect 23581 2261 23615 2295
rect 29929 2261 29963 2295
rect 36921 2261 36955 2295
<< metal1 >>
rect 1104 38650 37628 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 37628 38650
rect 1104 38576 37628 38598
rect 1762 38536 1768 38548
rect 1723 38508 1768 38536
rect 1762 38496 1768 38508
rect 1820 38496 1826 38548
rect 4706 38536 4712 38548
rect 4667 38508 4712 38536
rect 4706 38496 4712 38508
rect 4764 38496 4770 38548
rect 7650 38536 7656 38548
rect 7611 38508 7656 38536
rect 7650 38496 7656 38508
rect 7708 38496 7714 38548
rect 9861 38539 9919 38545
rect 9861 38505 9873 38539
rect 9907 38536 9919 38539
rect 10502 38536 10508 38548
rect 9907 38508 10508 38536
rect 9907 38505 9919 38508
rect 9861 38499 9919 38505
rect 10502 38496 10508 38508
rect 10560 38496 10566 38548
rect 11149 38539 11207 38545
rect 11149 38505 11161 38539
rect 11195 38536 11207 38539
rect 13078 38536 13084 38548
rect 11195 38508 13084 38536
rect 11195 38505 11207 38508
rect 11149 38499 11207 38505
rect 13078 38496 13084 38508
rect 13136 38496 13142 38548
rect 16298 38536 16304 38548
rect 16259 38508 16304 38536
rect 16298 38496 16304 38508
rect 16356 38496 16362 38548
rect 22278 38496 22284 38548
rect 22336 38536 22342 38548
rect 22373 38539 22431 38545
rect 22373 38536 22385 38539
rect 22336 38508 22385 38536
rect 22336 38496 22342 38508
rect 22373 38505 22385 38508
rect 22419 38505 22431 38539
rect 22373 38499 22431 38505
rect 25222 38496 25228 38548
rect 25280 38536 25286 38548
rect 25869 38539 25927 38545
rect 25869 38536 25881 38539
rect 25280 38508 25881 38536
rect 25280 38496 25286 38508
rect 25869 38505 25881 38508
rect 25915 38505 25927 38539
rect 25869 38499 25927 38505
rect 27709 38539 27767 38545
rect 27709 38505 27721 38539
rect 27755 38505 27767 38539
rect 27709 38499 27767 38505
rect 29917 38539 29975 38545
rect 29917 38505 29929 38539
rect 29963 38536 29975 38539
rect 30282 38536 30288 38548
rect 29963 38508 30288 38536
rect 29963 38505 29975 38508
rect 29917 38499 29975 38505
rect 12897 38471 12955 38477
rect 12897 38468 12909 38471
rect 6886 38440 12909 38468
rect 6886 38400 6914 38440
rect 12897 38437 12909 38440
rect 12943 38437 12955 38471
rect 12897 38431 12955 38437
rect 15289 38471 15347 38477
rect 15289 38437 15301 38471
rect 15335 38468 15347 38471
rect 19058 38468 19064 38480
rect 15335 38440 19064 38468
rect 15335 38437 15347 38440
rect 15289 38431 15347 38437
rect 19058 38428 19064 38440
rect 19116 38428 19122 38480
rect 27724 38468 27752 38499
rect 30282 38496 30288 38508
rect 30340 38496 30346 38548
rect 34054 38496 34060 38548
rect 34112 38536 34118 38548
rect 34149 38539 34207 38545
rect 34149 38536 34161 38539
rect 34112 38508 34161 38536
rect 34112 38496 34118 38508
rect 34149 38505 34161 38508
rect 34195 38505 34207 38539
rect 36906 38536 36912 38548
rect 36867 38508 36912 38536
rect 34149 38499 34207 38505
rect 36906 38496 36912 38508
rect 36964 38496 36970 38548
rect 23584 38440 27752 38468
rect 1964 38372 6914 38400
rect 18417 38403 18475 38409
rect 1964 38341 1992 38372
rect 18417 38369 18429 38403
rect 18463 38400 18475 38403
rect 18690 38400 18696 38412
rect 18463 38372 18696 38400
rect 18463 38369 18475 38372
rect 18417 38363 18475 38369
rect 18690 38360 18696 38372
rect 18748 38360 18754 38412
rect 19978 38400 19984 38412
rect 19939 38372 19984 38400
rect 19978 38360 19984 38372
rect 20036 38360 20042 38412
rect 20346 38360 20352 38412
rect 20404 38400 20410 38412
rect 20717 38403 20775 38409
rect 20717 38400 20729 38403
rect 20404 38372 20729 38400
rect 20404 38360 20410 38372
rect 20717 38369 20729 38372
rect 20763 38369 20775 38403
rect 20717 38363 20775 38369
rect 1949 38335 2007 38341
rect 1949 38301 1961 38335
rect 1995 38301 2007 38335
rect 1949 38295 2007 38301
rect 4798 38292 4804 38344
rect 4856 38332 4862 38344
rect 4893 38335 4951 38341
rect 4893 38332 4905 38335
rect 4856 38304 4905 38332
rect 4856 38292 4862 38304
rect 4893 38301 4905 38304
rect 4939 38301 4951 38335
rect 4893 38295 4951 38301
rect 7837 38335 7895 38341
rect 7837 38301 7849 38335
rect 7883 38332 7895 38335
rect 8110 38332 8116 38344
rect 7883 38304 8116 38332
rect 7883 38301 7895 38304
rect 7837 38295 7895 38301
rect 8110 38292 8116 38304
rect 8168 38292 8174 38344
rect 9677 38335 9735 38341
rect 9677 38301 9689 38335
rect 9723 38332 9735 38335
rect 10134 38332 10140 38344
rect 9723 38304 10140 38332
rect 9723 38301 9735 38304
rect 9677 38295 9735 38301
rect 10134 38292 10140 38304
rect 10192 38292 10198 38344
rect 10321 38335 10379 38341
rect 10321 38301 10333 38335
rect 10367 38332 10379 38335
rect 10410 38332 10416 38344
rect 10367 38304 10416 38332
rect 10367 38301 10379 38304
rect 10321 38295 10379 38301
rect 10410 38292 10416 38304
rect 10468 38292 10474 38344
rect 10965 38335 11023 38341
rect 10965 38332 10977 38335
rect 10520 38304 10977 38332
rect 10520 38205 10548 38304
rect 10965 38301 10977 38304
rect 11011 38301 11023 38335
rect 10965 38295 11023 38301
rect 12253 38335 12311 38341
rect 12253 38301 12265 38335
rect 12299 38301 12311 38335
rect 13078 38332 13084 38344
rect 13039 38304 13084 38332
rect 12253 38295 12311 38301
rect 12268 38264 12296 38295
rect 13078 38292 13084 38304
rect 13136 38292 13142 38344
rect 13541 38335 13599 38341
rect 13541 38301 13553 38335
rect 13587 38301 13599 38335
rect 14642 38332 14648 38344
rect 14603 38304 14648 38332
rect 13541 38295 13599 38301
rect 12618 38264 12624 38276
rect 12268 38236 12624 38264
rect 12618 38224 12624 38236
rect 12676 38264 12682 38276
rect 13556 38264 13584 38295
rect 14642 38292 14648 38304
rect 14700 38292 14706 38344
rect 15010 38292 15016 38344
rect 15068 38332 15074 38344
rect 15105 38335 15163 38341
rect 15105 38332 15117 38335
rect 15068 38304 15117 38332
rect 15068 38292 15074 38304
rect 15105 38301 15117 38304
rect 15151 38301 15163 38335
rect 15105 38295 15163 38301
rect 15746 38292 15752 38344
rect 15804 38332 15810 38344
rect 16117 38335 16175 38341
rect 16117 38332 16129 38335
rect 15804 38304 16129 38332
rect 15804 38292 15810 38304
rect 16117 38301 16129 38304
rect 16163 38301 16175 38335
rect 16117 38295 16175 38301
rect 17313 38335 17371 38341
rect 17313 38301 17325 38335
rect 17359 38332 17371 38335
rect 17359 38304 17816 38332
rect 17359 38301 17371 38304
rect 17313 38295 17371 38301
rect 12676 38236 13584 38264
rect 13633 38267 13691 38273
rect 12676 38224 12682 38236
rect 13633 38233 13645 38267
rect 13679 38264 13691 38267
rect 15194 38264 15200 38276
rect 13679 38236 15200 38264
rect 13679 38233 13691 38236
rect 13633 38227 13691 38233
rect 15194 38224 15200 38236
rect 15252 38224 15258 38276
rect 10505 38199 10563 38205
rect 10505 38165 10517 38199
rect 10551 38165 10563 38199
rect 12342 38196 12348 38208
rect 12303 38168 12348 38196
rect 10505 38159 10563 38165
rect 12342 38156 12348 38168
rect 12400 38156 12406 38208
rect 14090 38156 14096 38208
rect 14148 38196 14154 38208
rect 14461 38199 14519 38205
rect 14461 38196 14473 38199
rect 14148 38168 14473 38196
rect 14148 38156 14154 38168
rect 14461 38165 14473 38168
rect 14507 38165 14519 38199
rect 17126 38196 17132 38208
rect 17087 38168 17132 38196
rect 14461 38159 14519 38165
rect 17126 38156 17132 38168
rect 17184 38156 17190 38208
rect 17788 38205 17816 38304
rect 19518 38292 19524 38344
rect 19576 38332 19582 38344
rect 20993 38335 21051 38341
rect 20993 38332 21005 38335
rect 19576 38304 21005 38332
rect 19576 38292 19582 38304
rect 20993 38301 21005 38304
rect 21039 38301 21051 38335
rect 22554 38332 22560 38344
rect 22515 38304 22560 38332
rect 20993 38295 21051 38301
rect 18233 38267 18291 38273
rect 18233 38233 18245 38267
rect 18279 38264 18291 38267
rect 18598 38264 18604 38276
rect 18279 38236 18604 38264
rect 18279 38233 18291 38236
rect 18233 38227 18291 38233
rect 18598 38224 18604 38236
rect 18656 38264 18662 38276
rect 19797 38267 19855 38273
rect 19797 38264 19809 38267
rect 18656 38236 19809 38264
rect 18656 38224 18662 38236
rect 19797 38233 19809 38236
rect 19843 38264 19855 38267
rect 20901 38267 20959 38273
rect 20901 38264 20913 38267
rect 19843 38236 20913 38264
rect 19843 38233 19855 38236
rect 19797 38227 19855 38233
rect 20901 38233 20913 38236
rect 20947 38233 20959 38267
rect 21008 38264 21036 38295
rect 22554 38292 22560 38304
rect 22612 38292 22618 38344
rect 23017 38335 23075 38341
rect 23017 38301 23029 38335
rect 23063 38332 23075 38335
rect 23474 38332 23480 38344
rect 23063 38304 23480 38332
rect 23063 38301 23075 38304
rect 23017 38295 23075 38301
rect 23474 38292 23480 38304
rect 23532 38292 23538 38344
rect 23584 38276 23612 38440
rect 27724 38400 27752 38440
rect 28166 38428 28172 38480
rect 28224 38468 28230 38480
rect 30561 38471 30619 38477
rect 30561 38468 30573 38471
rect 28224 38440 30573 38468
rect 28224 38428 28230 38440
rect 30561 38437 30573 38440
rect 30607 38437 30619 38471
rect 30561 38431 30619 38437
rect 29546 38400 29552 38412
rect 27724 38372 29552 38400
rect 29546 38360 29552 38372
rect 29604 38360 29610 38412
rect 23658 38292 23664 38344
rect 23716 38332 23722 38344
rect 24762 38332 24768 38344
rect 23716 38304 23761 38332
rect 24723 38304 24768 38332
rect 23716 38292 23722 38304
rect 24762 38292 24768 38304
rect 24820 38292 24826 38344
rect 25406 38332 25412 38344
rect 25367 38304 25412 38332
rect 25406 38292 25412 38304
rect 25464 38292 25470 38344
rect 27985 38335 28043 38341
rect 27985 38301 27997 38335
rect 28031 38332 28043 38335
rect 28534 38332 28540 38344
rect 28031 38304 28540 38332
rect 28031 38301 28043 38304
rect 27985 38295 28043 38301
rect 28534 38292 28540 38304
rect 28592 38332 28598 38344
rect 28813 38335 28871 38341
rect 28813 38332 28825 38335
rect 28592 38304 28825 38332
rect 28592 38292 28598 38304
rect 28813 38301 28825 38304
rect 28859 38332 28871 38335
rect 31205 38335 31263 38341
rect 31205 38332 31217 38335
rect 28859 38304 29776 38332
rect 28859 38301 28871 38304
rect 28813 38295 28871 38301
rect 29748 38276 29776 38304
rect 30116 38304 31217 38332
rect 23566 38264 23572 38276
rect 21008 38236 23572 38264
rect 20901 38227 20959 38233
rect 23566 38224 23572 38236
rect 23624 38224 23630 38276
rect 29730 38264 29736 38276
rect 29643 38236 29736 38264
rect 29730 38224 29736 38236
rect 29788 38224 29794 38276
rect 30116 38208 30144 38304
rect 31205 38301 31217 38304
rect 31251 38301 31263 38335
rect 31386 38332 31392 38344
rect 31347 38304 31392 38332
rect 31205 38295 31263 38301
rect 31386 38292 31392 38304
rect 31444 38292 31450 38344
rect 32493 38335 32551 38341
rect 32493 38301 32505 38335
rect 32539 38332 32551 38335
rect 32953 38335 33011 38341
rect 32953 38332 32965 38335
rect 32539 38304 32965 38332
rect 32539 38301 32551 38304
rect 32493 38295 32551 38301
rect 32953 38301 32965 38304
rect 32999 38332 33011 38335
rect 33502 38332 33508 38344
rect 32999 38304 33508 38332
rect 32999 38301 33011 38304
rect 32953 38295 33011 38301
rect 33502 38292 33508 38304
rect 33560 38292 33566 38344
rect 34698 38292 34704 38344
rect 34756 38332 34762 38344
rect 36725 38335 36783 38341
rect 36725 38332 36737 38335
rect 34756 38304 36737 38332
rect 34756 38292 34762 38304
rect 36725 38301 36737 38304
rect 36771 38301 36783 38335
rect 36725 38295 36783 38301
rect 17773 38199 17831 38205
rect 17773 38165 17785 38199
rect 17819 38165 17831 38199
rect 18138 38196 18144 38208
rect 18099 38168 18144 38196
rect 17773 38159 17831 38165
rect 18138 38156 18144 38168
rect 18196 38156 18202 38208
rect 19426 38196 19432 38208
rect 19387 38168 19432 38196
rect 19426 38156 19432 38168
rect 19484 38156 19490 38208
rect 19886 38196 19892 38208
rect 19847 38168 19892 38196
rect 19886 38156 19892 38168
rect 19944 38156 19950 38208
rect 21358 38196 21364 38208
rect 21319 38168 21364 38196
rect 21358 38156 21364 38168
rect 21416 38156 21422 38208
rect 23106 38196 23112 38208
rect 23067 38168 23112 38196
rect 23106 38156 23112 38168
rect 23164 38156 23170 38208
rect 23750 38196 23756 38208
rect 23711 38168 23756 38196
rect 23750 38156 23756 38168
rect 23808 38156 23814 38208
rect 24486 38156 24492 38208
rect 24544 38196 24550 38208
rect 24581 38199 24639 38205
rect 24581 38196 24593 38199
rect 24544 38168 24593 38196
rect 24544 38156 24550 38168
rect 24581 38165 24593 38168
rect 24627 38165 24639 38199
rect 25222 38196 25228 38208
rect 25183 38168 25228 38196
rect 24581 38159 24639 38165
rect 25222 38156 25228 38168
rect 25280 38156 25286 38208
rect 27525 38199 27583 38205
rect 27525 38165 27537 38199
rect 27571 38196 27583 38199
rect 27706 38196 27712 38208
rect 27571 38168 27712 38196
rect 27571 38165 27583 38168
rect 27525 38159 27583 38165
rect 27706 38156 27712 38168
rect 27764 38156 27770 38208
rect 28718 38196 28724 38208
rect 28679 38168 28724 38196
rect 28718 38156 28724 38168
rect 28776 38156 28782 38208
rect 29914 38156 29920 38208
rect 29972 38205 29978 38208
rect 29972 38199 29991 38205
rect 29979 38165 29991 38199
rect 30098 38196 30104 38208
rect 30059 38168 30104 38196
rect 29972 38159 29991 38165
rect 29972 38156 29978 38159
rect 30098 38156 30104 38168
rect 30156 38156 30162 38208
rect 31297 38199 31355 38205
rect 31297 38165 31309 38199
rect 31343 38196 31355 38199
rect 31478 38196 31484 38208
rect 31343 38168 31484 38196
rect 31343 38165 31355 38168
rect 31297 38159 31355 38165
rect 31478 38156 31484 38168
rect 31536 38156 31542 38208
rect 32398 38196 32404 38208
rect 32359 38168 32404 38196
rect 32398 38156 32404 38168
rect 32456 38156 32462 38208
rect 33042 38196 33048 38208
rect 33003 38168 33048 38196
rect 33042 38156 33048 38168
rect 33100 38156 33106 38208
rect 1104 38106 37628 38128
rect 1104 38054 4874 38106
rect 4926 38054 4938 38106
rect 4990 38054 5002 38106
rect 5054 38054 5066 38106
rect 5118 38054 5130 38106
rect 5182 38054 35594 38106
rect 35646 38054 35658 38106
rect 35710 38054 35722 38106
rect 35774 38054 35786 38106
rect 35838 38054 35850 38106
rect 35902 38054 37628 38106
rect 1104 38032 37628 38054
rect 1578 37992 1584 38004
rect 1539 37964 1584 37992
rect 1578 37952 1584 37964
rect 1636 37952 1642 38004
rect 4798 37952 4804 38004
rect 4856 37992 4862 38004
rect 5077 37995 5135 38001
rect 5077 37992 5089 37995
rect 4856 37964 5089 37992
rect 4856 37952 4862 37964
rect 5077 37961 5089 37964
rect 5123 37961 5135 37995
rect 8110 37992 8116 38004
rect 8071 37964 8116 37992
rect 5077 37955 5135 37961
rect 8110 37952 8116 37964
rect 8168 37952 8174 38004
rect 10134 37992 10140 38004
rect 10095 37964 10140 37992
rect 10134 37952 10140 37964
rect 10192 37952 10198 38004
rect 12437 37995 12495 38001
rect 12437 37961 12449 37995
rect 12483 37961 12495 37995
rect 12437 37955 12495 37961
rect 12452 37924 12480 37955
rect 13078 37952 13084 38004
rect 13136 37992 13142 38004
rect 13909 37995 13967 38001
rect 13909 37992 13921 37995
rect 13136 37964 13921 37992
rect 13136 37952 13142 37964
rect 13909 37961 13921 37964
rect 13955 37961 13967 37995
rect 15746 37992 15752 38004
rect 15707 37964 15752 37992
rect 13909 37955 13967 37961
rect 15746 37952 15752 37964
rect 15804 37952 15810 38004
rect 18598 37992 18604 38004
rect 18559 37964 18604 37992
rect 18598 37952 18604 37964
rect 18656 37952 18662 38004
rect 19242 37992 19248 38004
rect 19203 37964 19248 37992
rect 19242 37952 19248 37964
rect 19300 37952 19306 38004
rect 21085 37995 21143 38001
rect 21085 37961 21097 37995
rect 21131 37992 21143 37995
rect 21131 37964 22324 37992
rect 21131 37961 21143 37964
rect 21085 37955 21143 37961
rect 17126 37924 17132 37936
rect 6886 37896 12480 37924
rect 14016 37896 14504 37924
rect 17087 37896 17132 37924
rect 1762 37856 1768 37868
rect 1723 37828 1768 37856
rect 1762 37816 1768 37828
rect 1820 37816 1826 37868
rect 5261 37859 5319 37865
rect 5261 37825 5273 37859
rect 5307 37856 5319 37859
rect 6886 37856 6914 37896
rect 8294 37856 8300 37868
rect 5307 37828 6914 37856
rect 8255 37828 8300 37856
rect 5307 37825 5319 37828
rect 5261 37819 5319 37825
rect 8294 37816 8300 37828
rect 8352 37816 8358 37868
rect 9582 37856 9588 37868
rect 9543 37828 9588 37856
rect 9582 37816 9588 37828
rect 9640 37816 9646 37868
rect 10318 37856 10324 37868
rect 10279 37828 10324 37856
rect 10318 37816 10324 37828
rect 10376 37816 10382 37868
rect 10778 37856 10784 37868
rect 10739 37828 10784 37856
rect 10778 37816 10784 37828
rect 10836 37816 10842 37868
rect 11606 37816 11612 37868
rect 11664 37856 11670 37868
rect 11793 37859 11851 37865
rect 11793 37856 11805 37859
rect 11664 37828 11805 37856
rect 11664 37816 11670 37828
rect 11793 37825 11805 37828
rect 11839 37825 11851 37859
rect 12802 37856 12808 37868
rect 12763 37828 12808 37856
rect 11793 37819 11851 37825
rect 12802 37816 12808 37828
rect 12860 37816 12866 37868
rect 12897 37859 12955 37865
rect 12897 37825 12909 37859
rect 12943 37856 12955 37859
rect 13446 37856 13452 37868
rect 12943 37828 13452 37856
rect 12943 37825 12955 37828
rect 12897 37819 12955 37825
rect 13446 37816 13452 37828
rect 13504 37816 13510 37868
rect 13081 37791 13139 37797
rect 13081 37757 13093 37791
rect 13127 37788 13139 37791
rect 14016 37788 14044 37896
rect 14274 37856 14280 37868
rect 14235 37828 14280 37856
rect 14274 37816 14280 37828
rect 14332 37816 14338 37868
rect 14476 37800 14504 37896
rect 17126 37884 17132 37896
rect 17184 37884 17190 37936
rect 19886 37884 19892 37936
rect 19944 37924 19950 37936
rect 20073 37927 20131 37933
rect 20073 37924 20085 37927
rect 19944 37896 20085 37924
rect 19944 37884 19950 37896
rect 20073 37893 20085 37896
rect 20119 37924 20131 37927
rect 22002 37924 22008 37936
rect 20119 37896 22008 37924
rect 20119 37893 20131 37896
rect 20073 37887 20131 37893
rect 22002 37884 22008 37896
rect 22060 37884 22066 37936
rect 22296 37933 22324 37964
rect 23750 37952 23756 38004
rect 23808 37992 23814 38004
rect 23808 37964 24716 37992
rect 23808 37952 23814 37964
rect 22281 37927 22339 37933
rect 22281 37893 22293 37927
rect 22327 37893 22339 37927
rect 22281 37887 22339 37893
rect 22738 37884 22744 37936
rect 22796 37884 22802 37936
rect 24486 37924 24492 37936
rect 24447 37896 24492 37924
rect 24486 37884 24492 37896
rect 24544 37884 24550 37936
rect 24688 37924 24716 37964
rect 29730 37952 29736 38004
rect 29788 37992 29794 38004
rect 30009 37995 30067 38001
rect 30009 37992 30021 37995
rect 29788 37964 30021 37992
rect 29788 37952 29794 37964
rect 30009 37961 30021 37964
rect 30055 37961 30067 37995
rect 33410 37992 33416 38004
rect 30009 37955 30067 37961
rect 31128 37964 33416 37992
rect 24688 37896 24978 37924
rect 15286 37816 15292 37868
rect 15344 37856 15350 37868
rect 15565 37859 15623 37865
rect 15565 37856 15577 37859
rect 15344 37828 15577 37856
rect 15344 37816 15350 37828
rect 15565 37825 15577 37828
rect 15611 37825 15623 37859
rect 15565 37819 15623 37825
rect 18230 37816 18236 37868
rect 18288 37816 18294 37868
rect 19058 37856 19064 37868
rect 19019 37828 19064 37856
rect 19058 37816 19064 37828
rect 19116 37816 19122 37868
rect 20901 37859 20959 37865
rect 20901 37825 20913 37859
rect 20947 37856 20959 37859
rect 21358 37856 21364 37868
rect 20947 37828 21364 37856
rect 20947 37825 20959 37828
rect 20901 37819 20959 37825
rect 21358 37816 21364 37828
rect 21416 37816 21422 37868
rect 24210 37856 24216 37868
rect 23492 37828 24216 37856
rect 14366 37788 14372 37800
rect 13127 37760 14044 37788
rect 14327 37760 14372 37788
rect 13127 37757 13139 37760
rect 13081 37751 13139 37757
rect 14366 37748 14372 37760
rect 14424 37748 14430 37800
rect 14458 37748 14464 37800
rect 14516 37788 14522 37800
rect 16850 37788 16856 37800
rect 14516 37760 14561 37788
rect 16811 37760 16856 37788
rect 14516 37748 14522 37760
rect 16850 37748 16856 37760
rect 16908 37748 16914 37800
rect 20162 37788 20168 37800
rect 20123 37760 20168 37788
rect 20162 37748 20168 37760
rect 20220 37748 20226 37800
rect 20346 37788 20352 37800
rect 20307 37760 20352 37788
rect 20346 37748 20352 37760
rect 20404 37748 20410 37800
rect 22005 37791 22063 37797
rect 22005 37757 22017 37791
rect 22051 37788 22063 37791
rect 23492 37788 23520 37828
rect 24210 37816 24216 37828
rect 24268 37816 24274 37868
rect 26418 37856 26424 37868
rect 26379 37828 26424 37856
rect 26418 37816 26424 37828
rect 26476 37816 26482 37868
rect 27154 37816 27160 37868
rect 27212 37856 27218 37868
rect 27249 37859 27307 37865
rect 27249 37856 27261 37859
rect 27212 37828 27261 37856
rect 27212 37816 27218 37828
rect 27249 37825 27261 37828
rect 27295 37856 27307 37859
rect 28074 37856 28080 37868
rect 27295 37828 28080 37856
rect 27295 37825 27307 37828
rect 27249 37819 27307 37825
rect 28074 37816 28080 37828
rect 28132 37816 28138 37868
rect 28169 37859 28227 37865
rect 28169 37825 28181 37859
rect 28215 37856 28227 37859
rect 29362 37856 29368 37868
rect 28215 37828 29368 37856
rect 28215 37825 28227 37828
rect 28169 37819 28227 37825
rect 22051 37760 23520 37788
rect 22051 37757 22063 37760
rect 22005 37751 22063 37757
rect 23566 37748 23572 37800
rect 23624 37788 23630 37800
rect 23753 37791 23811 37797
rect 23753 37788 23765 37791
rect 23624 37760 23765 37788
rect 23624 37748 23630 37760
rect 23753 37757 23765 37760
rect 23799 37757 23811 37791
rect 23753 37751 23811 37757
rect 11977 37723 12035 37729
rect 11977 37689 11989 37723
rect 12023 37720 12035 37723
rect 14734 37720 14740 37732
rect 12023 37692 14740 37720
rect 12023 37689 12035 37692
rect 11977 37683 12035 37689
rect 14734 37680 14740 37692
rect 14792 37680 14798 37732
rect 28184 37720 28212 37819
rect 29362 37816 29368 37828
rect 29420 37816 29426 37868
rect 29546 37856 29552 37868
rect 29507 37828 29552 37856
rect 29546 37816 29552 37828
rect 29604 37816 29610 37868
rect 27540 37692 28212 37720
rect 9398 37652 9404 37664
rect 9359 37624 9404 37652
rect 9398 37612 9404 37624
rect 9456 37612 9462 37664
rect 10962 37652 10968 37664
rect 10923 37624 10968 37652
rect 10962 37612 10968 37624
rect 11020 37612 11026 37664
rect 19610 37612 19616 37664
rect 19668 37652 19674 37664
rect 19705 37655 19763 37661
rect 19705 37652 19717 37655
rect 19668 37624 19717 37652
rect 19668 37612 19674 37624
rect 19705 37621 19717 37624
rect 19751 37621 19763 37655
rect 19705 37615 19763 37621
rect 25498 37612 25504 37664
rect 25556 37652 25562 37664
rect 25961 37655 26019 37661
rect 25961 37652 25973 37655
rect 25556 37624 25973 37652
rect 25556 37612 25562 37624
rect 25961 37621 25973 37624
rect 26007 37621 26019 37655
rect 26510 37652 26516 37664
rect 26471 37624 26516 37652
rect 25961 37615 26019 37621
rect 26510 37612 26516 37624
rect 26568 37612 26574 37664
rect 27540 37661 27568 37692
rect 27525 37655 27583 37661
rect 27525 37621 27537 37655
rect 27571 37621 27583 37655
rect 27525 37615 27583 37621
rect 27709 37655 27767 37661
rect 27709 37621 27721 37655
rect 27755 37652 27767 37655
rect 27982 37652 27988 37664
rect 27755 37624 27988 37652
rect 27755 37621 27767 37624
rect 27709 37615 27767 37621
rect 27982 37612 27988 37624
rect 28040 37612 28046 37664
rect 28074 37612 28080 37664
rect 28132 37652 28138 37664
rect 28261 37655 28319 37661
rect 28261 37652 28273 37655
rect 28132 37624 28273 37652
rect 28132 37612 28138 37624
rect 28261 37621 28273 37624
rect 28307 37621 28319 37655
rect 28626 37652 28632 37664
rect 28587 37624 28632 37652
rect 28261 37615 28319 37621
rect 28626 37612 28632 37624
rect 28684 37612 28690 37664
rect 29086 37652 29092 37664
rect 29047 37624 29092 37652
rect 29086 37612 29092 37624
rect 29144 37612 29150 37664
rect 29457 37655 29515 37661
rect 29457 37621 29469 37655
rect 29503 37652 29515 37655
rect 29748 37652 29776 37952
rect 31128 37924 31156 37964
rect 33410 37952 33416 37964
rect 33468 37952 33474 38004
rect 34698 37992 34704 38004
rect 34659 37964 34704 37992
rect 34698 37952 34704 37964
rect 34756 37952 34762 38004
rect 31478 37924 31484 37936
rect 31050 37896 31156 37924
rect 31439 37896 31484 37924
rect 31478 37884 31484 37896
rect 31536 37884 31542 37936
rect 33042 37884 33048 37936
rect 33100 37884 33106 37936
rect 34514 37856 34520 37868
rect 34475 37828 34520 37856
rect 34514 37816 34520 37828
rect 34572 37816 34578 37868
rect 31754 37748 31760 37800
rect 31812 37788 31818 37800
rect 33778 37788 33784 37800
rect 31812 37760 32812 37788
rect 33739 37760 33784 37788
rect 31812 37748 31818 37760
rect 29503 37624 29776 37652
rect 29503 37621 29515 37624
rect 29457 37615 29515 37621
rect 30282 37612 30288 37664
rect 30340 37652 30346 37664
rect 32309 37655 32367 37661
rect 32309 37652 32321 37655
rect 30340 37624 32321 37652
rect 30340 37612 30346 37624
rect 32309 37621 32321 37624
rect 32355 37621 32367 37655
rect 32784 37652 32812 37760
rect 33778 37748 33784 37760
rect 33836 37748 33842 37800
rect 34054 37788 34060 37800
rect 34015 37760 34060 37788
rect 34054 37748 34060 37760
rect 34112 37748 34118 37800
rect 34054 37652 34060 37664
rect 32784 37624 34060 37652
rect 32309 37615 32367 37621
rect 34054 37612 34060 37624
rect 34112 37612 34118 37664
rect 1104 37562 37628 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 37628 37562
rect 1104 37488 37628 37510
rect 13446 37448 13452 37460
rect 13407 37420 13452 37448
rect 13446 37408 13452 37420
rect 13504 37408 13510 37460
rect 14553 37451 14611 37457
rect 14553 37417 14565 37451
rect 14599 37448 14611 37451
rect 14642 37448 14648 37460
rect 14599 37420 14648 37448
rect 14599 37417 14611 37420
rect 14553 37411 14611 37417
rect 14642 37408 14648 37420
rect 14700 37408 14706 37460
rect 14734 37408 14740 37460
rect 14792 37448 14798 37460
rect 22554 37448 22560 37460
rect 14792 37420 22560 37448
rect 14792 37408 14798 37420
rect 22554 37408 22560 37420
rect 22612 37408 22618 37460
rect 24029 37451 24087 37457
rect 24029 37417 24041 37451
rect 24075 37448 24087 37451
rect 24762 37448 24768 37460
rect 24075 37420 24768 37448
rect 24075 37417 24087 37420
rect 24029 37411 24087 37417
rect 24762 37408 24768 37420
rect 24820 37408 24826 37460
rect 28074 37408 28080 37460
rect 28132 37448 28138 37460
rect 28261 37451 28319 37457
rect 28261 37448 28273 37451
rect 28132 37420 28273 37448
rect 28132 37408 28138 37420
rect 28261 37417 28273 37420
rect 28307 37417 28319 37451
rect 28261 37411 28319 37417
rect 30193 37451 30251 37457
rect 30193 37417 30205 37451
rect 30239 37448 30251 37451
rect 33778 37448 33784 37460
rect 30239 37420 33784 37448
rect 30239 37417 30251 37420
rect 30193 37411 30251 37417
rect 33778 37408 33784 37420
rect 33836 37408 33842 37460
rect 27706 37380 27712 37392
rect 27667 37352 27712 37380
rect 27706 37340 27712 37352
rect 27764 37380 27770 37392
rect 28810 37380 28816 37392
rect 27764 37352 28816 37380
rect 27764 37340 27770 37352
rect 28810 37340 28816 37352
rect 28868 37340 28874 37392
rect 9398 37312 9404 37324
rect 9359 37284 9404 37312
rect 9398 37272 9404 37284
rect 9456 37272 9462 37324
rect 13814 37272 13820 37324
rect 13872 37312 13878 37324
rect 15102 37312 15108 37324
rect 13872 37284 15108 37312
rect 13872 37272 13878 37284
rect 15102 37272 15108 37284
rect 15160 37272 15166 37324
rect 18325 37315 18383 37321
rect 18325 37281 18337 37315
rect 18371 37312 18383 37315
rect 18690 37312 18696 37324
rect 18371 37284 18696 37312
rect 18371 37281 18383 37284
rect 18325 37275 18383 37281
rect 18690 37272 18696 37284
rect 18748 37272 18754 37324
rect 23477 37315 23535 37321
rect 23477 37281 23489 37315
rect 23523 37312 23535 37315
rect 23566 37312 23572 37324
rect 23523 37284 23572 37312
rect 23523 37281 23535 37284
rect 23477 37275 23535 37281
rect 23566 37272 23572 37284
rect 23624 37272 23630 37324
rect 24210 37272 24216 37324
rect 24268 37312 24274 37324
rect 24854 37312 24860 37324
rect 24268 37284 24860 37312
rect 24268 37272 24274 37284
rect 24854 37272 24860 37284
rect 24912 37312 24918 37324
rect 24949 37315 25007 37321
rect 24949 37312 24961 37315
rect 24912 37284 24961 37312
rect 24912 37272 24918 37284
rect 24949 37281 24961 37284
rect 24995 37281 25007 37315
rect 25222 37312 25228 37324
rect 25183 37284 25228 37312
rect 24949 37275 25007 37281
rect 25222 37272 25228 37284
rect 25280 37272 25286 37324
rect 27982 37272 27988 37324
rect 28040 37312 28046 37324
rect 30006 37312 30012 37324
rect 28040 37284 28856 37312
rect 29967 37284 30012 37312
rect 28040 37272 28046 37284
rect 8110 37204 8116 37256
rect 8168 37244 8174 37256
rect 8389 37247 8447 37253
rect 8389 37244 8401 37247
rect 8168 37216 8401 37244
rect 8168 37204 8174 37216
rect 8389 37213 8401 37216
rect 8435 37213 8447 37247
rect 8389 37207 8447 37213
rect 9125 37247 9183 37253
rect 9125 37213 9137 37247
rect 9171 37213 9183 37247
rect 9125 37207 9183 37213
rect 11701 37247 11759 37253
rect 11701 37213 11713 37247
rect 11747 37213 11759 37247
rect 11701 37207 11759 37213
rect 8202 37136 8208 37188
rect 8260 37176 8266 37188
rect 9140 37176 9168 37207
rect 8260 37148 9168 37176
rect 9232 37148 9890 37176
rect 8260 37136 8266 37148
rect 8481 37111 8539 37117
rect 8481 37077 8493 37111
rect 8527 37108 8539 37111
rect 9232 37108 9260 37148
rect 10870 37108 10876 37120
rect 8527 37080 9260 37108
rect 10831 37080 10876 37108
rect 8527 37077 8539 37080
rect 8481 37071 8539 37077
rect 10870 37068 10876 37080
rect 10928 37068 10934 37120
rect 11716 37108 11744 37207
rect 14366 37204 14372 37256
rect 14424 37244 14430 37256
rect 14918 37244 14924 37256
rect 14424 37216 14924 37244
rect 14424 37204 14430 37216
rect 14918 37204 14924 37216
rect 14976 37204 14982 37256
rect 15749 37247 15807 37253
rect 15749 37213 15761 37247
rect 15795 37213 15807 37247
rect 15749 37207 15807 37213
rect 18509 37247 18567 37253
rect 18509 37213 18521 37247
rect 18555 37244 18567 37247
rect 19426 37244 19432 37256
rect 18555 37216 19432 37244
rect 18555 37213 18567 37216
rect 18509 37207 18567 37213
rect 11974 37176 11980 37188
rect 11935 37148 11980 37176
rect 11974 37136 11980 37148
rect 12032 37136 12038 37188
rect 12360 37148 12466 37176
rect 12360 37120 12388 37148
rect 12250 37108 12256 37120
rect 11716 37080 12256 37108
rect 12250 37068 12256 37080
rect 12308 37068 12314 37120
rect 12342 37068 12348 37120
rect 12400 37068 12406 37120
rect 15013 37111 15071 37117
rect 15013 37077 15025 37111
rect 15059 37108 15071 37111
rect 15378 37108 15384 37120
rect 15059 37080 15384 37108
rect 15059 37077 15071 37080
rect 15013 37071 15071 37077
rect 15378 37068 15384 37080
rect 15436 37068 15442 37120
rect 15764 37108 15792 37207
rect 19426 37204 19432 37216
rect 19484 37204 19490 37256
rect 19610 37244 19616 37256
rect 19571 37216 19616 37244
rect 19610 37204 19616 37216
rect 19668 37204 19674 37256
rect 20254 37244 20260 37256
rect 20215 37216 20260 37244
rect 20254 37204 20260 37216
rect 20312 37204 20318 37256
rect 22741 37247 22799 37253
rect 22741 37213 22753 37247
rect 22787 37244 22799 37247
rect 23014 37244 23020 37256
rect 22787 37216 23020 37244
rect 22787 37213 22799 37216
rect 22741 37207 22799 37213
rect 23014 37204 23020 37216
rect 23072 37204 23078 37256
rect 27893 37247 27951 37253
rect 27893 37213 27905 37247
rect 27939 37244 27951 37247
rect 28626 37244 28632 37256
rect 27939 37216 28632 37244
rect 27939 37213 27951 37216
rect 27893 37207 27951 37213
rect 28626 37204 28632 37216
rect 28684 37244 28690 37256
rect 28721 37247 28779 37253
rect 28721 37244 28733 37247
rect 28684 37216 28733 37244
rect 28684 37204 28690 37216
rect 28721 37213 28733 37216
rect 28767 37213 28779 37247
rect 28828 37244 28856 37284
rect 30006 37272 30012 37284
rect 30064 37272 30070 37324
rect 31294 37312 31300 37324
rect 31036 37284 31300 37312
rect 29181 37247 29239 37253
rect 29181 37244 29193 37247
rect 28828 37216 29193 37244
rect 28721 37207 28779 37213
rect 29181 37213 29193 37216
rect 29227 37213 29239 37247
rect 29181 37207 29239 37213
rect 29270 37204 29276 37256
rect 29328 37244 29334 37256
rect 31036 37253 31064 37284
rect 31294 37272 31300 37284
rect 31352 37312 31358 37324
rect 31754 37312 31760 37324
rect 31352 37284 31760 37312
rect 31352 37272 31358 37284
rect 31754 37272 31760 37284
rect 31812 37272 31818 37324
rect 29917 37247 29975 37253
rect 29917 37244 29929 37247
rect 29328 37216 29929 37244
rect 29328 37204 29334 37216
rect 29917 37213 29929 37216
rect 29963 37213 29975 37247
rect 29917 37207 29975 37213
rect 31021 37247 31079 37253
rect 31021 37213 31033 37247
rect 31067 37213 31079 37247
rect 31021 37207 31079 37213
rect 32398 37204 32404 37256
rect 32456 37204 32462 37256
rect 33410 37244 33416 37256
rect 33371 37216 33416 37244
rect 33410 37204 33416 37216
rect 33468 37204 33474 37256
rect 33502 37204 33508 37256
rect 33560 37244 33566 37256
rect 33560 37216 33605 37244
rect 33560 37204 33566 37216
rect 16022 37176 16028 37188
rect 15983 37148 16028 37176
rect 16022 37136 16028 37148
rect 16080 37136 16086 37188
rect 17034 37136 17040 37188
rect 17092 37136 17098 37188
rect 18322 37136 18328 37188
rect 18380 37176 18386 37188
rect 18417 37179 18475 37185
rect 18417 37176 18429 37179
rect 18380 37148 18429 37176
rect 18380 37136 18386 37148
rect 18417 37145 18429 37148
rect 18463 37176 18475 37179
rect 20162 37176 20168 37188
rect 18463 37148 20168 37176
rect 18463 37145 18475 37148
rect 18417 37139 18475 37145
rect 20162 37136 20168 37148
rect 20220 37136 20226 37188
rect 20533 37179 20591 37185
rect 20533 37145 20545 37179
rect 20579 37145 20591 37179
rect 20533 37139 20591 37145
rect 16850 37108 16856 37120
rect 15764 37080 16856 37108
rect 16850 37068 16856 37080
rect 16908 37108 16914 37120
rect 17310 37108 17316 37120
rect 16908 37080 17316 37108
rect 16908 37068 16914 37080
rect 17310 37068 17316 37080
rect 17368 37068 17374 37120
rect 17497 37111 17555 37117
rect 17497 37077 17509 37111
rect 17543 37108 17555 37111
rect 17954 37108 17960 37120
rect 17543 37080 17960 37108
rect 17543 37077 17555 37080
rect 17497 37071 17555 37077
rect 17954 37068 17960 37080
rect 18012 37108 18018 37120
rect 18598 37108 18604 37120
rect 18012 37080 18604 37108
rect 18012 37068 18018 37080
rect 18598 37068 18604 37080
rect 18656 37068 18662 37120
rect 18877 37111 18935 37117
rect 18877 37077 18889 37111
rect 18923 37108 18935 37111
rect 19702 37108 19708 37120
rect 18923 37080 19708 37108
rect 18923 37077 18935 37080
rect 18877 37071 18935 37077
rect 19702 37068 19708 37080
rect 19760 37068 19766 37120
rect 19797 37111 19855 37117
rect 19797 37077 19809 37111
rect 19843 37108 19855 37111
rect 20548 37108 20576 37139
rect 21266 37136 21272 37188
rect 21324 37136 21330 37188
rect 23569 37179 23627 37185
rect 23569 37145 23581 37179
rect 23615 37176 23627 37179
rect 25498 37176 25504 37188
rect 23615 37148 25504 37176
rect 23615 37145 23627 37148
rect 23569 37139 23627 37145
rect 25498 37136 25504 37148
rect 25556 37136 25562 37188
rect 26510 37176 26516 37188
rect 26450 37148 26516 37176
rect 26510 37136 26516 37148
rect 26568 37136 26574 37188
rect 27982 37176 27988 37188
rect 27943 37148 27988 37176
rect 27982 37136 27988 37148
rect 28040 37136 28046 37188
rect 28077 37179 28135 37185
rect 28077 37145 28089 37179
rect 28123 37176 28135 37179
rect 29086 37176 29092 37188
rect 28123 37148 29092 37176
rect 28123 37145 28135 37148
rect 28077 37139 28135 37145
rect 29086 37136 29092 37148
rect 29144 37136 29150 37188
rect 30374 37136 30380 37188
rect 30432 37176 30438 37188
rect 31297 37179 31355 37185
rect 31297 37176 31309 37179
rect 30432 37148 31309 37176
rect 30432 37136 30438 37148
rect 31297 37145 31309 37148
rect 31343 37145 31355 37179
rect 31297 37139 31355 37145
rect 22002 37108 22008 37120
rect 19843 37080 20576 37108
rect 21963 37080 22008 37108
rect 19843 37077 19855 37080
rect 19797 37071 19855 37077
rect 22002 37068 22008 37080
rect 22060 37068 22066 37120
rect 22370 37068 22376 37120
rect 22428 37108 22434 37120
rect 22557 37111 22615 37117
rect 22557 37108 22569 37111
rect 22428 37080 22569 37108
rect 22428 37068 22434 37080
rect 22557 37077 22569 37080
rect 22603 37077 22615 37111
rect 22557 37071 22615 37077
rect 23658 37068 23664 37120
rect 23716 37108 23722 37120
rect 26694 37108 26700 37120
rect 23716 37080 23761 37108
rect 26655 37080 26700 37108
rect 23716 37068 23722 37080
rect 26694 37068 26700 37080
rect 26752 37068 26758 37120
rect 28810 37108 28816 37120
rect 28771 37080 28816 37108
rect 28810 37068 28816 37080
rect 28868 37068 28874 37120
rect 28902 37068 28908 37120
rect 28960 37108 28966 37120
rect 28960 37080 29005 37108
rect 28960 37068 28966 37080
rect 29362 37068 29368 37120
rect 29420 37108 29426 37120
rect 29822 37108 29828 37120
rect 29420 37080 29828 37108
rect 29420 37068 29426 37080
rect 29822 37068 29828 37080
rect 29880 37108 29886 37120
rect 32769 37111 32827 37117
rect 32769 37108 32781 37111
rect 29880 37080 32781 37108
rect 29880 37068 29886 37080
rect 32769 37077 32781 37080
rect 32815 37077 32827 37111
rect 32769 37071 32827 37077
rect 1104 37018 37628 37040
rect 1104 36966 4874 37018
rect 4926 36966 4938 37018
rect 4990 36966 5002 37018
rect 5054 36966 5066 37018
rect 5118 36966 5130 37018
rect 5182 36966 35594 37018
rect 35646 36966 35658 37018
rect 35710 36966 35722 37018
rect 35774 36966 35786 37018
rect 35838 36966 35850 37018
rect 35902 36966 37628 37018
rect 1104 36944 37628 36966
rect 8294 36864 8300 36916
rect 8352 36904 8358 36916
rect 9769 36907 9827 36913
rect 9769 36904 9781 36907
rect 8352 36876 9781 36904
rect 8352 36864 8358 36876
rect 9769 36873 9781 36876
rect 9815 36873 9827 36907
rect 9769 36867 9827 36873
rect 11149 36907 11207 36913
rect 11149 36873 11161 36907
rect 11195 36904 11207 36907
rect 11974 36904 11980 36916
rect 11195 36876 11980 36904
rect 11195 36873 11207 36876
rect 11149 36867 11207 36873
rect 11974 36864 11980 36876
rect 12032 36864 12038 36916
rect 12621 36907 12679 36913
rect 12621 36873 12633 36907
rect 12667 36873 12679 36907
rect 12621 36867 12679 36873
rect 12989 36907 13047 36913
rect 12989 36873 13001 36907
rect 13035 36904 13047 36907
rect 13446 36904 13452 36916
rect 13035 36876 13452 36904
rect 13035 36873 13047 36876
rect 12989 36867 13047 36873
rect 10137 36839 10195 36845
rect 10137 36805 10149 36839
rect 10183 36836 10195 36839
rect 10226 36836 10232 36848
rect 10183 36808 10232 36836
rect 10183 36805 10195 36808
rect 10137 36799 10195 36805
rect 10226 36796 10232 36808
rect 10284 36796 10290 36848
rect 12636 36836 12664 36867
rect 13446 36864 13452 36876
rect 13504 36864 13510 36916
rect 14918 36864 14924 36916
rect 14976 36904 14982 36916
rect 15565 36907 15623 36913
rect 15565 36904 15577 36907
rect 14976 36876 15577 36904
rect 14976 36864 14982 36876
rect 15565 36873 15577 36876
rect 15611 36873 15623 36907
rect 15565 36867 15623 36873
rect 16022 36864 16028 36916
rect 16080 36904 16086 36916
rect 16117 36907 16175 36913
rect 16117 36904 16129 36907
rect 16080 36876 16129 36904
rect 16080 36864 16086 36876
rect 16117 36873 16129 36876
rect 16163 36873 16175 36907
rect 16945 36907 17003 36913
rect 16945 36904 16957 36907
rect 16117 36867 16175 36873
rect 16546 36876 16957 36904
rect 13814 36836 13820 36848
rect 10980 36808 12664 36836
rect 13280 36808 13820 36836
rect 9217 36771 9275 36777
rect 9217 36737 9229 36771
rect 9263 36768 9275 36771
rect 9398 36768 9404 36780
rect 9263 36740 9404 36768
rect 9263 36737 9275 36740
rect 9217 36731 9275 36737
rect 9398 36728 9404 36740
rect 9456 36728 9462 36780
rect 10870 36768 10876 36780
rect 10244 36740 10876 36768
rect 9950 36660 9956 36712
rect 10008 36700 10014 36712
rect 10244 36709 10272 36740
rect 10870 36728 10876 36740
rect 10928 36728 10934 36780
rect 10980 36777 11008 36808
rect 10965 36771 11023 36777
rect 10965 36737 10977 36771
rect 11011 36737 11023 36771
rect 10965 36731 11023 36737
rect 11238 36728 11244 36780
rect 11296 36768 11302 36780
rect 12069 36771 12127 36777
rect 12069 36768 12081 36771
rect 11296 36740 12081 36768
rect 11296 36728 11302 36740
rect 12069 36737 12081 36740
rect 12115 36737 12127 36771
rect 12069 36731 12127 36737
rect 10229 36703 10287 36709
rect 10229 36700 10241 36703
rect 10008 36672 10241 36700
rect 10008 36660 10014 36672
rect 10229 36669 10241 36672
rect 10275 36669 10287 36703
rect 10229 36663 10287 36669
rect 10413 36703 10471 36709
rect 10413 36669 10425 36703
rect 10459 36700 10471 36703
rect 10594 36700 10600 36712
rect 10459 36672 10600 36700
rect 10459 36669 10471 36672
rect 10413 36663 10471 36669
rect 10594 36660 10600 36672
rect 10652 36660 10658 36712
rect 12618 36700 12624 36712
rect 10704 36672 12624 36700
rect 8110 36592 8116 36644
rect 8168 36632 8174 36644
rect 10704 36632 10732 36672
rect 12618 36660 12624 36672
rect 12676 36660 12682 36712
rect 13078 36700 13084 36712
rect 13039 36672 13084 36700
rect 13078 36660 13084 36672
rect 13136 36660 13142 36712
rect 13280 36709 13308 36808
rect 13814 36796 13820 36808
rect 13872 36796 13878 36848
rect 14090 36836 14096 36848
rect 14051 36808 14096 36836
rect 14090 36796 14096 36808
rect 14148 36796 14154 36848
rect 15194 36728 15200 36780
rect 15252 36728 15258 36780
rect 16301 36771 16359 36777
rect 16301 36737 16313 36771
rect 16347 36768 16359 36771
rect 16546 36768 16574 36876
rect 16945 36873 16957 36876
rect 16991 36873 17003 36907
rect 16945 36867 17003 36873
rect 17313 36907 17371 36913
rect 17313 36873 17325 36907
rect 17359 36904 17371 36907
rect 17954 36904 17960 36916
rect 17359 36876 17960 36904
rect 17359 36873 17371 36876
rect 17313 36867 17371 36873
rect 17954 36864 17960 36876
rect 18012 36864 18018 36916
rect 18141 36907 18199 36913
rect 18141 36873 18153 36907
rect 18187 36904 18199 36907
rect 18322 36904 18328 36916
rect 18187 36876 18328 36904
rect 18187 36873 18199 36876
rect 18141 36867 18199 36873
rect 18322 36864 18328 36876
rect 18380 36864 18386 36916
rect 20349 36907 20407 36913
rect 20349 36904 20361 36907
rect 19628 36876 20361 36904
rect 19150 36796 19156 36848
rect 19208 36796 19214 36848
rect 19628 36845 19656 36876
rect 20349 36873 20361 36876
rect 20395 36873 20407 36907
rect 20349 36867 20407 36873
rect 21266 36864 21272 36916
rect 21324 36904 21330 36916
rect 21361 36907 21419 36913
rect 21361 36904 21373 36907
rect 21324 36876 21373 36904
rect 21324 36864 21330 36876
rect 21361 36873 21373 36876
rect 21407 36873 21419 36907
rect 21361 36867 21419 36873
rect 23658 36864 23664 36916
rect 23716 36904 23722 36916
rect 24305 36907 24363 36913
rect 24305 36904 24317 36907
rect 23716 36876 24317 36904
rect 23716 36864 23722 36876
rect 24305 36873 24317 36876
rect 24351 36873 24363 36907
rect 24305 36867 24363 36873
rect 24394 36864 24400 36916
rect 24452 36904 24458 36916
rect 29003 36907 29061 36913
rect 24452 36876 28028 36904
rect 24452 36864 24458 36876
rect 28000 36848 28028 36876
rect 29003 36873 29015 36907
rect 29049 36904 29061 36907
rect 31386 36904 31392 36916
rect 29049 36876 31392 36904
rect 29049 36873 29061 36876
rect 29003 36867 29061 36873
rect 31386 36864 31392 36876
rect 31444 36864 31450 36916
rect 19613 36839 19671 36845
rect 19613 36805 19625 36839
rect 19659 36805 19671 36839
rect 19613 36799 19671 36805
rect 19702 36796 19708 36848
rect 19760 36836 19766 36848
rect 22370 36836 22376 36848
rect 19760 36808 20576 36836
rect 22331 36808 22376 36836
rect 19760 36796 19766 36808
rect 16347 36740 16574 36768
rect 17405 36771 17463 36777
rect 16347 36737 16359 36740
rect 16301 36731 16359 36737
rect 17405 36737 17417 36771
rect 17451 36768 17463 36771
rect 18322 36768 18328 36780
rect 17451 36740 18328 36768
rect 17451 36737 17463 36740
rect 17405 36731 17463 36737
rect 18322 36728 18328 36740
rect 18380 36728 18386 36780
rect 20548 36777 20576 36808
rect 22370 36796 22376 36808
rect 22428 36796 22434 36848
rect 23106 36796 23112 36848
rect 23164 36796 23170 36848
rect 24765 36839 24823 36845
rect 24765 36805 24777 36839
rect 24811 36836 24823 36839
rect 25869 36839 25927 36845
rect 25869 36836 25881 36839
rect 24811 36808 25881 36836
rect 24811 36805 24823 36808
rect 24765 36799 24823 36805
rect 25869 36805 25881 36808
rect 25915 36836 25927 36839
rect 26694 36836 26700 36848
rect 25915 36808 26700 36836
rect 25915 36805 25927 36808
rect 25869 36799 25927 36805
rect 26694 36796 26700 36808
rect 26752 36836 26758 36848
rect 27982 36836 27988 36848
rect 26752 36808 27200 36836
rect 27895 36808 27988 36836
rect 26752 36796 26758 36808
rect 20533 36771 20591 36777
rect 20533 36737 20545 36771
rect 20579 36737 20591 36771
rect 21266 36768 21272 36780
rect 21227 36740 21272 36768
rect 20533 36731 20591 36737
rect 21266 36728 21272 36740
rect 21324 36728 21330 36780
rect 24673 36771 24731 36777
rect 24673 36768 24685 36771
rect 23860 36740 24685 36768
rect 13265 36703 13323 36709
rect 13265 36669 13277 36703
rect 13311 36669 13323 36703
rect 13814 36700 13820 36712
rect 13775 36672 13820 36700
rect 13265 36663 13323 36669
rect 13814 36660 13820 36672
rect 13872 36660 13878 36712
rect 15102 36660 15108 36712
rect 15160 36700 15166 36712
rect 17126 36700 17132 36712
rect 15160 36672 17132 36700
rect 15160 36660 15166 36672
rect 17126 36660 17132 36672
rect 17184 36700 17190 36712
rect 17497 36703 17555 36709
rect 17497 36700 17509 36703
rect 17184 36672 17509 36700
rect 17184 36660 17190 36672
rect 17497 36669 17509 36672
rect 17543 36669 17555 36703
rect 17497 36663 17555 36669
rect 19889 36703 19947 36709
rect 19889 36669 19901 36703
rect 19935 36700 19947 36703
rect 20254 36700 20260 36712
rect 19935 36672 20260 36700
rect 19935 36669 19947 36672
rect 19889 36663 19947 36669
rect 8168 36604 10732 36632
rect 8168 36592 8174 36604
rect 9122 36564 9128 36576
rect 9083 36536 9128 36564
rect 9122 36524 9128 36536
rect 9180 36524 9186 36576
rect 11977 36567 12035 36573
rect 11977 36533 11989 36567
rect 12023 36564 12035 36567
rect 12066 36564 12072 36576
rect 12023 36536 12072 36564
rect 12023 36533 12035 36536
rect 11977 36527 12035 36533
rect 12066 36524 12072 36536
rect 12124 36524 12130 36576
rect 19426 36524 19432 36576
rect 19484 36564 19490 36576
rect 19904 36564 19932 36663
rect 20254 36660 20260 36672
rect 20312 36660 20318 36712
rect 22094 36700 22100 36712
rect 22055 36672 22100 36700
rect 22094 36660 22100 36672
rect 22152 36660 22158 36712
rect 19484 36536 19932 36564
rect 19484 36524 19490 36536
rect 23474 36524 23480 36576
rect 23532 36564 23538 36576
rect 23860 36573 23888 36740
rect 24673 36737 24685 36740
rect 24719 36737 24731 36771
rect 24673 36731 24731 36737
rect 25498 36728 25504 36780
rect 25556 36768 25562 36780
rect 25961 36771 26019 36777
rect 25961 36768 25973 36771
rect 25556 36740 25973 36768
rect 25556 36728 25562 36740
rect 25961 36737 25973 36740
rect 26007 36768 26019 36771
rect 26142 36768 26148 36780
rect 26007 36740 26148 36768
rect 26007 36737 26019 36740
rect 25961 36731 26019 36737
rect 26142 36728 26148 36740
rect 26200 36728 26206 36780
rect 27172 36777 27200 36808
rect 27982 36796 27988 36808
rect 28040 36796 28046 36848
rect 28534 36796 28540 36848
rect 28592 36836 28598 36848
rect 28905 36839 28963 36845
rect 28905 36836 28917 36839
rect 28592 36808 28917 36836
rect 28592 36796 28598 36808
rect 28905 36805 28917 36808
rect 28951 36805 28963 36839
rect 28905 36799 28963 36805
rect 29089 36839 29147 36845
rect 29089 36805 29101 36839
rect 29135 36836 29147 36839
rect 34054 36836 34060 36848
rect 29135 36808 30328 36836
rect 34015 36808 34060 36836
rect 29135 36805 29147 36808
rect 29089 36799 29147 36805
rect 27157 36771 27215 36777
rect 27157 36737 27169 36771
rect 27203 36737 27215 36771
rect 27157 36731 27215 36737
rect 24857 36703 24915 36709
rect 24857 36669 24869 36703
rect 24903 36669 24915 36703
rect 24857 36663 24915 36669
rect 23845 36567 23903 36573
rect 23845 36564 23857 36567
rect 23532 36536 23857 36564
rect 23532 36524 23538 36536
rect 23845 36533 23857 36536
rect 23891 36533 23903 36567
rect 23845 36527 23903 36533
rect 24026 36524 24032 36576
rect 24084 36564 24090 36576
rect 24872 36564 24900 36663
rect 24946 36660 24952 36712
rect 25004 36700 25010 36712
rect 26053 36703 26111 36709
rect 26053 36700 26065 36703
rect 25004 36672 26065 36700
rect 25004 36660 25010 36672
rect 26053 36669 26065 36672
rect 26099 36669 26111 36703
rect 26053 36663 26111 36669
rect 25406 36592 25412 36644
rect 25464 36632 25470 36644
rect 25501 36635 25559 36641
rect 25501 36632 25513 36635
rect 25464 36604 25513 36632
rect 25464 36592 25470 36604
rect 25501 36601 25513 36604
rect 25547 36601 25559 36635
rect 25501 36595 25559 36601
rect 28353 36635 28411 36641
rect 28353 36601 28365 36635
rect 28399 36632 28411 36635
rect 29104 36632 29132 36799
rect 30300 36780 30328 36808
rect 34054 36796 34060 36808
rect 34112 36796 34118 36848
rect 29181 36771 29239 36777
rect 29181 36737 29193 36771
rect 29227 36768 29239 36771
rect 29227 36740 29776 36768
rect 29227 36737 29239 36740
rect 29181 36731 29239 36737
rect 28399 36604 29132 36632
rect 29748 36632 29776 36740
rect 29822 36728 29828 36780
rect 29880 36768 29886 36780
rect 29880 36740 29925 36768
rect 29880 36728 29886 36740
rect 30282 36728 30288 36780
rect 30340 36768 30346 36780
rect 30837 36771 30895 36777
rect 30837 36768 30849 36771
rect 30340 36740 30849 36768
rect 30340 36728 30346 36740
rect 30837 36737 30849 36740
rect 30883 36737 30895 36771
rect 30837 36731 30895 36737
rect 32309 36771 32367 36777
rect 32309 36737 32321 36771
rect 32355 36768 32367 36771
rect 33594 36768 33600 36780
rect 32355 36740 33600 36768
rect 32355 36737 32367 36740
rect 32309 36731 32367 36737
rect 33594 36728 33600 36740
rect 33652 36728 33658 36780
rect 29917 36703 29975 36709
rect 29917 36669 29929 36703
rect 29963 36700 29975 36703
rect 30098 36700 30104 36712
rect 29963 36672 30104 36700
rect 29963 36669 29975 36672
rect 29917 36663 29975 36669
rect 30098 36660 30104 36672
rect 30156 36660 30162 36712
rect 30193 36703 30251 36709
rect 30193 36669 30205 36703
rect 30239 36700 30251 36703
rect 30374 36700 30380 36712
rect 30239 36672 30380 36700
rect 30239 36669 30251 36672
rect 30193 36663 30251 36669
rect 30374 36660 30380 36672
rect 30432 36660 30438 36712
rect 30006 36632 30012 36644
rect 29748 36604 30012 36632
rect 28399 36601 28411 36604
rect 28353 36595 28411 36601
rect 30006 36592 30012 36604
rect 30064 36592 30070 36644
rect 27246 36564 27252 36576
rect 24084 36536 24900 36564
rect 27207 36536 27252 36564
rect 24084 36524 24090 36536
rect 27246 36524 27252 36536
rect 27304 36524 27310 36576
rect 28166 36524 28172 36576
rect 28224 36564 28230 36576
rect 28445 36567 28503 36573
rect 28445 36564 28457 36567
rect 28224 36536 28457 36564
rect 28224 36524 28230 36536
rect 28445 36533 28457 36536
rect 28491 36533 28503 36567
rect 28445 36527 28503 36533
rect 29086 36524 29092 36576
rect 29144 36564 29150 36576
rect 30745 36567 30803 36573
rect 30745 36564 30757 36567
rect 29144 36536 30757 36564
rect 29144 36524 29150 36536
rect 30745 36533 30757 36536
rect 30791 36533 30803 36567
rect 30745 36527 30803 36533
rect 1104 36474 37628 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 37628 36474
rect 1104 36400 37628 36422
rect 9582 36360 9588 36372
rect 9543 36332 9588 36360
rect 9582 36320 9588 36332
rect 9640 36320 9646 36372
rect 11238 36360 11244 36372
rect 9692 36332 11244 36360
rect 9398 36252 9404 36304
rect 9456 36292 9462 36304
rect 9692 36292 9720 36332
rect 11238 36320 11244 36332
rect 11296 36320 11302 36372
rect 16945 36363 17003 36369
rect 16945 36329 16957 36363
rect 16991 36360 17003 36363
rect 17034 36360 17040 36372
rect 16991 36332 17040 36360
rect 16991 36329 17003 36332
rect 16945 36323 17003 36329
rect 17034 36320 17040 36332
rect 17092 36320 17098 36372
rect 18138 36360 18144 36372
rect 18099 36332 18144 36360
rect 18138 36320 18144 36332
rect 18196 36320 18202 36372
rect 21913 36363 21971 36369
rect 21913 36329 21925 36363
rect 21959 36360 21971 36363
rect 22738 36360 22744 36372
rect 21959 36332 22744 36360
rect 21959 36329 21971 36332
rect 21913 36323 21971 36329
rect 22738 36320 22744 36332
rect 22796 36320 22802 36372
rect 23014 36360 23020 36372
rect 22975 36332 23020 36360
rect 23014 36320 23020 36332
rect 23072 36320 23078 36372
rect 27154 36360 27160 36372
rect 25240 36332 27160 36360
rect 9456 36264 9720 36292
rect 9456 36252 9462 36264
rect 12250 36252 12256 36304
rect 12308 36292 12314 36304
rect 13814 36292 13820 36304
rect 12308 36264 13820 36292
rect 12308 36252 12314 36264
rect 13814 36252 13820 36264
rect 13872 36252 13878 36304
rect 17589 36295 17647 36301
rect 17589 36261 17601 36295
rect 17635 36292 17647 36295
rect 18230 36292 18236 36304
rect 17635 36264 18236 36292
rect 17635 36261 17647 36264
rect 17589 36255 17647 36261
rect 18230 36252 18236 36264
rect 18288 36252 18294 36304
rect 18598 36252 18604 36304
rect 18656 36292 18662 36304
rect 25240 36292 25268 36332
rect 27154 36320 27160 36332
rect 27212 36320 27218 36372
rect 30101 36363 30159 36369
rect 30101 36329 30113 36363
rect 30147 36360 30159 36363
rect 30282 36360 30288 36372
rect 30147 36332 30288 36360
rect 30147 36329 30159 36332
rect 30101 36323 30159 36329
rect 30282 36320 30288 36332
rect 30340 36320 30346 36372
rect 31202 36320 31208 36372
rect 31260 36360 31266 36372
rect 33045 36363 33103 36369
rect 33045 36360 33057 36363
rect 31260 36332 33057 36360
rect 31260 36320 31266 36332
rect 33045 36329 33057 36332
rect 33091 36329 33103 36363
rect 33045 36323 33103 36329
rect 18656 36264 25268 36292
rect 25317 36295 25375 36301
rect 18656 36252 18662 36264
rect 25317 36261 25329 36295
rect 25363 36261 25375 36295
rect 25317 36255 25375 36261
rect 27985 36295 28043 36301
rect 27985 36261 27997 36295
rect 28031 36261 28043 36295
rect 27985 36255 28043 36261
rect 28721 36295 28779 36301
rect 28721 36261 28733 36295
rect 28767 36292 28779 36295
rect 28994 36292 29000 36304
rect 28767 36264 29000 36292
rect 28767 36261 28779 36264
rect 28721 36255 28779 36261
rect 8018 36184 8024 36236
rect 8076 36224 8082 36236
rect 8481 36227 8539 36233
rect 8481 36224 8493 36227
rect 8076 36196 8493 36224
rect 8076 36184 8082 36196
rect 8481 36193 8493 36196
rect 8527 36224 8539 36227
rect 10229 36227 10287 36233
rect 10229 36224 10241 36227
rect 8527 36196 10241 36224
rect 8527 36193 8539 36196
rect 8481 36187 8539 36193
rect 10229 36193 10241 36196
rect 10275 36224 10287 36227
rect 12434 36224 12440 36236
rect 10275 36196 12440 36224
rect 10275 36193 10287 36196
rect 10229 36187 10287 36193
rect 12434 36184 12440 36196
rect 12492 36184 12498 36236
rect 13446 36224 13452 36236
rect 13407 36196 13452 36224
rect 13446 36184 13452 36196
rect 13504 36184 13510 36236
rect 13633 36227 13691 36233
rect 13633 36193 13645 36227
rect 13679 36224 13691 36227
rect 14921 36227 14979 36233
rect 14921 36224 14933 36227
rect 13679 36196 14933 36224
rect 13679 36193 13691 36196
rect 13633 36187 13691 36193
rect 14921 36193 14933 36196
rect 14967 36224 14979 36227
rect 16022 36224 16028 36236
rect 14967 36196 16028 36224
rect 14967 36193 14979 36196
rect 14921 36187 14979 36193
rect 16022 36184 16028 36196
rect 16080 36224 16086 36236
rect 18785 36227 18843 36233
rect 18785 36224 18797 36227
rect 16080 36196 18797 36224
rect 16080 36184 16086 36196
rect 18785 36193 18797 36196
rect 18831 36224 18843 36227
rect 19702 36224 19708 36236
rect 18831 36196 19708 36224
rect 18831 36193 18843 36196
rect 18785 36187 18843 36193
rect 19702 36184 19708 36196
rect 19760 36224 19766 36236
rect 19889 36227 19947 36233
rect 19889 36224 19901 36227
rect 19760 36196 19901 36224
rect 19760 36184 19766 36196
rect 19889 36193 19901 36196
rect 19935 36224 19947 36227
rect 19978 36224 19984 36236
rect 19935 36196 19984 36224
rect 19935 36193 19947 36196
rect 19889 36187 19947 36193
rect 19978 36184 19984 36196
rect 20036 36184 20042 36236
rect 23474 36224 23480 36236
rect 23435 36196 23480 36224
rect 23474 36184 23480 36196
rect 23532 36184 23538 36236
rect 23566 36184 23572 36236
rect 23624 36224 23630 36236
rect 24765 36227 24823 36233
rect 23624 36196 23669 36224
rect 23624 36184 23630 36196
rect 24765 36193 24777 36227
rect 24811 36224 24823 36227
rect 24946 36224 24952 36236
rect 24811 36196 24952 36224
rect 24811 36193 24823 36196
rect 24765 36187 24823 36193
rect 24946 36184 24952 36196
rect 25004 36184 25010 36236
rect 7098 36116 7104 36168
rect 7156 36156 7162 36168
rect 7193 36159 7251 36165
rect 7193 36156 7205 36159
rect 7156 36128 7205 36156
rect 7156 36116 7162 36128
rect 7193 36125 7205 36128
rect 7239 36156 7251 36159
rect 8110 36156 8116 36168
rect 7239 36128 8116 36156
rect 7239 36125 7251 36128
rect 7193 36119 7251 36125
rect 8110 36116 8116 36128
rect 8168 36116 8174 36168
rect 9950 36156 9956 36168
rect 9911 36128 9956 36156
rect 9950 36116 9956 36128
rect 10008 36116 10014 36168
rect 10410 36116 10416 36168
rect 10468 36156 10474 36168
rect 10781 36159 10839 36165
rect 10781 36156 10793 36159
rect 10468 36128 10793 36156
rect 10468 36116 10474 36128
rect 10781 36125 10793 36128
rect 10827 36125 10839 36159
rect 10781 36119 10839 36125
rect 13078 36116 13084 36168
rect 13136 36156 13142 36168
rect 15197 36159 15255 36165
rect 15197 36156 15209 36159
rect 13136 36128 15209 36156
rect 13136 36116 13142 36128
rect 15197 36125 15209 36128
rect 15243 36125 15255 36159
rect 17034 36156 17040 36168
rect 16995 36128 17040 36156
rect 15197 36119 15255 36125
rect 17034 36116 17040 36128
rect 17092 36116 17098 36168
rect 17678 36156 17684 36168
rect 17639 36128 17684 36156
rect 17678 36116 17684 36128
rect 17736 36116 17742 36168
rect 17954 36116 17960 36168
rect 18012 36156 18018 36168
rect 18322 36156 18328 36168
rect 18012 36128 18328 36156
rect 18012 36116 18018 36128
rect 18322 36116 18328 36128
rect 18380 36156 18386 36168
rect 18509 36159 18567 36165
rect 18509 36156 18521 36159
rect 18380 36128 18521 36156
rect 18380 36116 18386 36128
rect 18509 36125 18521 36128
rect 18555 36125 18567 36159
rect 18509 36119 18567 36125
rect 18601 36159 18659 36165
rect 18601 36125 18613 36159
rect 18647 36156 18659 36159
rect 19518 36156 19524 36168
rect 18647 36128 19524 36156
rect 18647 36125 18659 36128
rect 18601 36119 18659 36125
rect 19518 36116 19524 36128
rect 19576 36116 19582 36168
rect 20073 36159 20131 36165
rect 20073 36125 20085 36159
rect 20119 36156 20131 36159
rect 20162 36156 20168 36168
rect 20119 36128 20168 36156
rect 20119 36125 20131 36128
rect 20073 36119 20131 36125
rect 20162 36116 20168 36128
rect 20220 36116 20226 36168
rect 21821 36159 21879 36165
rect 21821 36125 21833 36159
rect 21867 36125 21879 36159
rect 23492 36156 23520 36184
rect 24857 36159 24915 36165
rect 24857 36156 24869 36159
rect 23492 36128 24869 36156
rect 21821 36119 21879 36125
rect 24857 36125 24869 36128
rect 24903 36125 24915 36159
rect 25332 36156 25360 36255
rect 27614 36184 27620 36236
rect 27672 36224 27678 36236
rect 28000 36224 28028 36255
rect 28994 36252 29000 36264
rect 29052 36252 29058 36304
rect 31294 36224 31300 36236
rect 27672 36196 30604 36224
rect 31255 36196 31300 36224
rect 27672 36184 27678 36196
rect 30576 36168 30604 36196
rect 31294 36184 31300 36196
rect 31352 36224 31358 36236
rect 32306 36224 32312 36236
rect 31352 36196 32312 36224
rect 31352 36184 31358 36196
rect 32306 36184 32312 36196
rect 32364 36184 32370 36236
rect 25961 36159 26019 36165
rect 25961 36156 25973 36159
rect 25332 36128 25973 36156
rect 24857 36119 24915 36125
rect 25961 36125 25973 36128
rect 26007 36125 26019 36159
rect 26418 36156 26424 36168
rect 26331 36128 26424 36156
rect 25961 36119 26019 36125
rect 10962 36048 10968 36100
rect 11020 36088 11026 36100
rect 11057 36091 11115 36097
rect 11057 36088 11069 36091
rect 11020 36060 11069 36088
rect 11020 36048 11026 36060
rect 11057 36057 11069 36060
rect 11103 36057 11115 36091
rect 11057 36051 11115 36057
rect 12066 36048 12072 36100
rect 12124 36048 12130 36100
rect 13357 36091 13415 36097
rect 13357 36088 13369 36091
rect 12544 36060 13369 36088
rect 7285 36023 7343 36029
rect 7285 35989 7297 36023
rect 7331 36020 7343 36023
rect 7374 36020 7380 36032
rect 7331 35992 7380 36020
rect 7331 35989 7343 35992
rect 7285 35983 7343 35989
rect 7374 35980 7380 35992
rect 7432 35980 7438 36032
rect 7466 35980 7472 36032
rect 7524 36020 7530 36032
rect 7837 36023 7895 36029
rect 7837 36020 7849 36023
rect 7524 35992 7849 36020
rect 7524 35980 7530 35992
rect 7837 35989 7849 35992
rect 7883 35989 7895 36023
rect 7837 35983 7895 35989
rect 8110 35980 8116 36032
rect 8168 36020 8174 36032
rect 8205 36023 8263 36029
rect 8205 36020 8217 36023
rect 8168 35992 8217 36020
rect 8168 35980 8174 35992
rect 8205 35989 8217 35992
rect 8251 35989 8263 36023
rect 8205 35983 8263 35989
rect 8294 35980 8300 36032
rect 8352 36020 8358 36032
rect 10045 36023 10103 36029
rect 8352 35992 8397 36020
rect 8352 35980 8358 35992
rect 10045 35989 10057 36023
rect 10091 36020 10103 36023
rect 10686 36020 10692 36032
rect 10091 35992 10692 36020
rect 10091 35989 10103 35992
rect 10045 35983 10103 35989
rect 10686 35980 10692 35992
rect 10744 36020 10750 36032
rect 12544 36029 12572 36060
rect 13357 36057 13369 36060
rect 13403 36057 13415 36091
rect 13357 36051 13415 36057
rect 14918 36048 14924 36100
rect 14976 36088 14982 36100
rect 15105 36091 15163 36097
rect 15105 36088 15117 36091
rect 14976 36060 15117 36088
rect 14976 36048 14982 36060
rect 15105 36057 15117 36060
rect 15151 36057 15163 36091
rect 15105 36051 15163 36057
rect 17310 36048 17316 36100
rect 17368 36088 17374 36100
rect 19426 36088 19432 36100
rect 17368 36060 19432 36088
rect 17368 36048 17374 36060
rect 19426 36048 19432 36060
rect 19484 36048 19490 36100
rect 21266 36048 21272 36100
rect 21324 36088 21330 36100
rect 21836 36088 21864 36119
rect 26418 36116 26424 36128
rect 26476 36116 26482 36168
rect 27982 36116 27988 36168
rect 28040 36156 28046 36168
rect 30193 36159 30251 36165
rect 30193 36156 30205 36159
rect 28040 36128 30205 36156
rect 28040 36116 28046 36128
rect 30193 36125 30205 36128
rect 30239 36125 30251 36159
rect 30193 36119 30251 36125
rect 30558 36116 30564 36168
rect 30616 36156 30622 36168
rect 30653 36159 30711 36165
rect 30653 36156 30665 36159
rect 30616 36128 30665 36156
rect 30616 36116 30622 36128
rect 30653 36125 30665 36128
rect 30699 36125 30711 36159
rect 30834 36156 30840 36168
rect 30795 36128 30840 36156
rect 30653 36119 30711 36125
rect 30834 36116 30840 36128
rect 30892 36116 30898 36168
rect 33502 36116 33508 36168
rect 33560 36156 33566 36168
rect 33689 36159 33747 36165
rect 33689 36156 33701 36159
rect 33560 36128 33701 36156
rect 33560 36116 33566 36128
rect 33689 36125 33701 36128
rect 33735 36125 33747 36159
rect 33689 36119 33747 36125
rect 26436 36088 26464 36116
rect 21324 36060 26464 36088
rect 21324 36048 21330 36060
rect 26970 36048 26976 36100
rect 27028 36088 27034 36100
rect 27617 36091 27675 36097
rect 27617 36088 27629 36091
rect 27028 36060 27629 36088
rect 27028 36048 27034 36060
rect 27617 36057 27629 36060
rect 27663 36057 27675 36091
rect 27617 36051 27675 36057
rect 28442 36048 28448 36100
rect 28500 36088 28506 36100
rect 28997 36091 29055 36097
rect 28997 36088 29009 36091
rect 28500 36060 29009 36088
rect 28500 36048 28506 36060
rect 28997 36057 29009 36060
rect 29043 36057 29055 36091
rect 28997 36051 29055 36057
rect 30282 36048 30288 36100
rect 30340 36088 30346 36100
rect 31573 36091 31631 36097
rect 31573 36088 31585 36091
rect 30340 36060 31585 36088
rect 30340 36048 30346 36060
rect 31573 36057 31585 36060
rect 31619 36057 31631 36091
rect 33042 36088 33048 36100
rect 32798 36060 33048 36088
rect 31573 36051 31631 36057
rect 33042 36048 33048 36060
rect 33100 36048 33106 36100
rect 12529 36023 12587 36029
rect 12529 36020 12541 36023
rect 10744 35992 12541 36020
rect 10744 35980 10750 35992
rect 12529 35989 12541 35992
rect 12575 35989 12587 36023
rect 12986 36020 12992 36032
rect 12947 35992 12992 36020
rect 12529 35983 12587 35989
rect 12986 35980 12992 35992
rect 13044 35980 13050 36032
rect 15562 36020 15568 36032
rect 15523 35992 15568 36020
rect 15562 35980 15568 35992
rect 15620 35980 15626 36032
rect 19978 36020 19984 36032
rect 19939 35992 19984 36020
rect 19978 35980 19984 35992
rect 20036 35980 20042 36032
rect 20438 36020 20444 36032
rect 20399 35992 20444 36020
rect 20438 35980 20444 35992
rect 20496 35980 20502 36032
rect 23382 36020 23388 36032
rect 23343 35992 23388 36020
rect 23382 35980 23388 35992
rect 23440 35980 23446 36032
rect 24946 36020 24952 36032
rect 24907 35992 24952 36020
rect 24946 35980 24952 35992
rect 25004 35980 25010 36032
rect 25130 35980 25136 36032
rect 25188 36020 25194 36032
rect 25777 36023 25835 36029
rect 25777 36020 25789 36023
rect 25188 35992 25789 36020
rect 25188 35980 25194 35992
rect 25777 35989 25789 35992
rect 25823 35989 25835 36023
rect 26510 36020 26516 36032
rect 26471 35992 26516 36020
rect 25777 35983 25835 35989
rect 26510 35980 26516 35992
rect 26568 35980 26574 36032
rect 28077 36023 28135 36029
rect 28077 35989 28089 36023
rect 28123 36020 28135 36023
rect 28258 36020 28264 36032
rect 28123 35992 28264 36020
rect 28123 35989 28135 35992
rect 28077 35983 28135 35989
rect 28258 35980 28264 35992
rect 28316 35980 28322 36032
rect 28534 36020 28540 36032
rect 28495 35992 28540 36020
rect 28534 35980 28540 35992
rect 28592 35980 28598 36032
rect 29730 36020 29736 36032
rect 29691 35992 29736 36020
rect 29730 35980 29736 35992
rect 29788 35980 29794 36032
rect 30745 36023 30803 36029
rect 30745 35989 30757 36023
rect 30791 36020 30803 36023
rect 31662 36020 31668 36032
rect 30791 35992 31668 36020
rect 30791 35989 30803 35992
rect 30745 35983 30803 35989
rect 31662 35980 31668 35992
rect 31720 35980 31726 36032
rect 33597 36023 33655 36029
rect 33597 35989 33609 36023
rect 33643 36020 33655 36023
rect 33686 36020 33692 36032
rect 33643 35992 33692 36020
rect 33643 35989 33655 35992
rect 33597 35983 33655 35989
rect 33686 35980 33692 35992
rect 33744 35980 33750 36032
rect 1104 35930 37628 35952
rect 1104 35878 4874 35930
rect 4926 35878 4938 35930
rect 4990 35878 5002 35930
rect 5054 35878 5066 35930
rect 5118 35878 5130 35930
rect 5182 35878 35594 35930
rect 35646 35878 35658 35930
rect 35710 35878 35722 35930
rect 35774 35878 35786 35930
rect 35838 35878 35850 35930
rect 35902 35878 37628 35930
rect 1104 35856 37628 35878
rect 10686 35816 10692 35828
rect 10647 35788 10692 35816
rect 10686 35776 10692 35788
rect 10744 35776 10750 35828
rect 10778 35776 10784 35828
rect 10836 35816 10842 35828
rect 11149 35819 11207 35825
rect 11149 35816 11161 35819
rect 10836 35788 11161 35816
rect 10836 35776 10842 35788
rect 11149 35785 11161 35788
rect 11195 35785 11207 35819
rect 11149 35779 11207 35785
rect 12986 35776 12992 35828
rect 13044 35816 13050 35828
rect 13265 35819 13323 35825
rect 13265 35816 13277 35819
rect 13044 35788 13277 35816
rect 13044 35776 13050 35788
rect 13265 35785 13277 35788
rect 13311 35785 13323 35819
rect 13265 35779 13323 35785
rect 13633 35819 13691 35825
rect 13633 35785 13645 35819
rect 13679 35785 13691 35819
rect 13633 35779 13691 35785
rect 15289 35819 15347 35825
rect 15289 35785 15301 35819
rect 15335 35816 15347 35819
rect 15562 35816 15568 35828
rect 15335 35788 15568 35816
rect 15335 35785 15347 35788
rect 15289 35779 15347 35785
rect 7466 35748 7472 35760
rect 6886 35720 7472 35748
rect 6549 35683 6607 35689
rect 6549 35649 6561 35683
rect 6595 35680 6607 35683
rect 6886 35680 6914 35720
rect 7466 35708 7472 35720
rect 7524 35708 7530 35760
rect 8202 35748 8208 35760
rect 7852 35720 8208 35748
rect 7190 35680 7196 35692
rect 6595 35652 6914 35680
rect 7151 35652 7196 35680
rect 6595 35649 6607 35652
rect 6549 35643 6607 35649
rect 7190 35640 7196 35652
rect 7248 35640 7254 35692
rect 7852 35689 7880 35720
rect 8202 35708 8208 35720
rect 8260 35708 8266 35760
rect 9122 35708 9128 35760
rect 9180 35708 9186 35760
rect 9950 35708 9956 35760
rect 10008 35748 10014 35760
rect 12161 35751 12219 35757
rect 12161 35748 12173 35751
rect 10008 35720 12173 35748
rect 10008 35708 10014 35720
rect 12161 35717 12173 35720
rect 12207 35717 12219 35751
rect 13648 35748 13676 35779
rect 15562 35776 15568 35788
rect 15620 35776 15626 35828
rect 19150 35816 19156 35828
rect 19111 35788 19156 35816
rect 19150 35776 19156 35788
rect 19208 35776 19214 35828
rect 20165 35819 20223 35825
rect 20165 35785 20177 35819
rect 20211 35816 20223 35819
rect 20438 35816 20444 35828
rect 20211 35788 20444 35816
rect 20211 35785 20223 35788
rect 20165 35779 20223 35785
rect 20438 35776 20444 35788
rect 20496 35776 20502 35828
rect 23382 35776 23388 35828
rect 23440 35816 23446 35828
rect 23477 35819 23535 35825
rect 23477 35816 23489 35819
rect 23440 35788 23489 35816
rect 23440 35776 23446 35788
rect 23477 35785 23489 35788
rect 23523 35785 23535 35819
rect 23477 35779 23535 35785
rect 23937 35819 23995 35825
rect 23937 35785 23949 35819
rect 23983 35816 23995 35819
rect 24946 35816 24952 35828
rect 23983 35788 24952 35816
rect 23983 35785 23995 35788
rect 23937 35779 23995 35785
rect 24946 35776 24952 35788
rect 25004 35816 25010 35828
rect 26605 35819 26663 35825
rect 26605 35816 26617 35819
rect 25004 35788 26617 35816
rect 25004 35776 25010 35788
rect 26605 35785 26617 35788
rect 26651 35785 26663 35819
rect 26605 35779 26663 35785
rect 27985 35819 28043 35825
rect 27985 35785 27997 35819
rect 28031 35816 28043 35819
rect 34057 35819 34115 35825
rect 34057 35816 34069 35819
rect 28031 35788 28856 35816
rect 28031 35785 28043 35788
rect 27985 35779 28043 35785
rect 13648 35720 16344 35748
rect 12161 35711 12219 35717
rect 7837 35683 7895 35689
rect 7837 35649 7849 35683
rect 7883 35649 7895 35683
rect 7837 35643 7895 35649
rect 10781 35683 10839 35689
rect 10781 35649 10793 35683
rect 10827 35649 10839 35683
rect 10781 35643 10839 35649
rect 12069 35683 12127 35689
rect 12069 35649 12081 35683
rect 12115 35649 12127 35683
rect 14274 35680 14280 35692
rect 14235 35652 14280 35680
rect 12069 35643 12127 35649
rect 8113 35615 8171 35621
rect 8113 35612 8125 35615
rect 7392 35584 8125 35612
rect 7392 35553 7420 35584
rect 8113 35581 8125 35584
rect 8159 35581 8171 35615
rect 8113 35575 8171 35581
rect 10597 35615 10655 35621
rect 10597 35581 10609 35615
rect 10643 35612 10655 35615
rect 10686 35612 10692 35624
rect 10643 35584 10692 35612
rect 10643 35581 10655 35584
rect 10597 35575 10655 35581
rect 10686 35572 10692 35584
rect 10744 35572 10750 35624
rect 7377 35547 7435 35553
rect 7377 35513 7389 35547
rect 7423 35513 7435 35547
rect 10796 35544 10824 35643
rect 11701 35547 11759 35553
rect 11701 35544 11713 35547
rect 10796 35516 11713 35544
rect 7377 35507 7435 35513
rect 11701 35513 11713 35516
rect 11747 35513 11759 35547
rect 11701 35507 11759 35513
rect 6730 35476 6736 35488
rect 6691 35448 6736 35476
rect 6730 35436 6736 35448
rect 6788 35436 6794 35488
rect 8294 35436 8300 35488
rect 8352 35476 8358 35488
rect 9582 35476 9588 35488
rect 8352 35448 9588 35476
rect 8352 35436 8358 35448
rect 9582 35436 9588 35448
rect 9640 35476 9646 35488
rect 12084 35476 12112 35643
rect 14274 35640 14280 35652
rect 14332 35640 14338 35692
rect 15378 35680 15384 35692
rect 15291 35652 15384 35680
rect 15378 35640 15384 35652
rect 15436 35680 15442 35692
rect 15930 35680 15936 35692
rect 15436 35652 15936 35680
rect 15436 35640 15442 35652
rect 15930 35640 15936 35652
rect 15988 35640 15994 35692
rect 16316 35689 16344 35720
rect 17678 35708 17684 35760
rect 17736 35748 17742 35760
rect 17736 35720 19288 35748
rect 17736 35708 17742 35720
rect 19260 35692 19288 35720
rect 19886 35708 19892 35760
rect 19944 35748 19950 35760
rect 20073 35751 20131 35757
rect 20073 35748 20085 35751
rect 19944 35720 20085 35748
rect 19944 35708 19950 35720
rect 20073 35717 20085 35720
rect 20119 35748 20131 35751
rect 22370 35748 22376 35760
rect 20119 35720 22376 35748
rect 20119 35717 20131 35720
rect 20073 35711 20131 35717
rect 22370 35708 22376 35720
rect 22428 35748 22434 35760
rect 23845 35751 23903 35757
rect 23845 35748 23857 35751
rect 22428 35720 23857 35748
rect 22428 35708 22434 35720
rect 23845 35717 23857 35720
rect 23891 35717 23903 35751
rect 25130 35748 25136 35760
rect 25091 35720 25136 35748
rect 23845 35711 23903 35717
rect 25130 35708 25136 35720
rect 25188 35708 25194 35760
rect 26510 35748 26516 35760
rect 26358 35720 26516 35748
rect 26510 35708 26516 35720
rect 26568 35708 26574 35760
rect 26620 35748 26648 35779
rect 28828 35760 28856 35788
rect 29932 35788 34069 35816
rect 29932 35760 29960 35788
rect 34057 35785 34069 35788
rect 34103 35785 34115 35819
rect 34057 35779 34115 35785
rect 28442 35748 28448 35760
rect 26620 35720 28448 35748
rect 28442 35708 28448 35720
rect 28500 35708 28506 35760
rect 28810 35748 28816 35760
rect 28723 35720 28816 35748
rect 28810 35708 28816 35720
rect 28868 35708 28874 35760
rect 28994 35708 29000 35760
rect 29052 35748 29058 35760
rect 29825 35751 29883 35757
rect 29825 35748 29837 35751
rect 29052 35720 29837 35748
rect 29052 35708 29058 35720
rect 29825 35717 29837 35720
rect 29871 35748 29883 35751
rect 29914 35748 29920 35760
rect 29871 35720 29920 35748
rect 29871 35717 29883 35720
rect 29825 35711 29883 35717
rect 29914 35708 29920 35720
rect 29972 35708 29978 35760
rect 30041 35751 30099 35757
rect 30041 35717 30053 35751
rect 30087 35748 30099 35751
rect 30374 35748 30380 35760
rect 30087 35720 30380 35748
rect 30087 35717 30099 35720
rect 30041 35711 30099 35717
rect 30374 35708 30380 35720
rect 30432 35708 30438 35760
rect 31202 35748 31208 35760
rect 30484 35720 31208 35748
rect 16301 35683 16359 35689
rect 16301 35649 16313 35683
rect 16347 35649 16359 35683
rect 17862 35680 17868 35692
rect 17823 35652 17868 35680
rect 16301 35643 16359 35649
rect 17862 35640 17868 35652
rect 17920 35640 17926 35692
rect 19242 35680 19248 35692
rect 19203 35652 19248 35680
rect 19242 35640 19248 35652
rect 19300 35640 19306 35692
rect 21177 35683 21235 35689
rect 21177 35680 21189 35683
rect 20548 35652 21189 35680
rect 12158 35572 12164 35624
rect 12216 35612 12222 35624
rect 12253 35615 12311 35621
rect 12253 35612 12265 35615
rect 12216 35584 12265 35612
rect 12216 35572 12222 35584
rect 12253 35581 12265 35584
rect 12299 35581 12311 35615
rect 12253 35575 12311 35581
rect 12989 35615 13047 35621
rect 12989 35581 13001 35615
rect 13035 35581 13047 35615
rect 13170 35612 13176 35624
rect 13131 35584 13176 35612
rect 12989 35575 13047 35581
rect 13004 35544 13032 35575
rect 13170 35572 13176 35584
rect 13228 35572 13234 35624
rect 13906 35612 13912 35624
rect 13280 35584 13912 35612
rect 13280 35544 13308 35584
rect 13906 35572 13912 35584
rect 13964 35612 13970 35624
rect 15102 35612 15108 35624
rect 13964 35584 15108 35612
rect 13964 35572 13970 35584
rect 15102 35572 15108 35584
rect 15160 35612 15166 35624
rect 15473 35615 15531 35621
rect 15473 35612 15485 35615
rect 15160 35584 15485 35612
rect 15160 35572 15166 35584
rect 15473 35581 15485 35584
rect 15519 35581 15531 35615
rect 17954 35612 17960 35624
rect 17915 35584 17960 35612
rect 15473 35575 15531 35581
rect 17954 35572 17960 35584
rect 18012 35572 18018 35624
rect 18141 35615 18199 35621
rect 18141 35581 18153 35615
rect 18187 35612 18199 35615
rect 18690 35612 18696 35624
rect 18187 35584 18696 35612
rect 18187 35581 18199 35584
rect 18141 35575 18199 35581
rect 18690 35572 18696 35584
rect 18748 35612 18754 35624
rect 19518 35612 19524 35624
rect 18748 35584 19524 35612
rect 18748 35572 18754 35584
rect 19518 35572 19524 35584
rect 19576 35612 19582 35624
rect 19889 35615 19947 35621
rect 19889 35612 19901 35615
rect 19576 35584 19901 35612
rect 19576 35572 19582 35584
rect 19889 35581 19901 35584
rect 19935 35581 19947 35615
rect 19889 35575 19947 35581
rect 13004 35516 13308 35544
rect 13538 35504 13544 35556
rect 13596 35544 13602 35556
rect 20548 35553 20576 35652
rect 21177 35649 21189 35652
rect 21223 35649 21235 35683
rect 21177 35643 21235 35649
rect 21358 35640 21364 35692
rect 21416 35680 21422 35692
rect 22189 35683 22247 35689
rect 22189 35680 22201 35683
rect 21416 35652 22201 35680
rect 21416 35640 21422 35652
rect 22189 35649 22201 35652
rect 22235 35649 22247 35683
rect 22189 35643 22247 35649
rect 22925 35683 22983 35689
rect 22925 35649 22937 35683
rect 22971 35680 22983 35683
rect 23290 35680 23296 35692
rect 22971 35652 23296 35680
rect 22971 35649 22983 35652
rect 22925 35643 22983 35649
rect 22204 35612 22232 35643
rect 23290 35640 23296 35652
rect 23348 35640 23354 35692
rect 24854 35680 24860 35692
rect 24815 35652 24860 35680
rect 24854 35640 24860 35652
rect 24912 35640 24918 35692
rect 28074 35680 28080 35692
rect 28035 35652 28080 35680
rect 28074 35640 28080 35652
rect 28132 35640 28138 35692
rect 28169 35683 28227 35689
rect 28169 35649 28181 35683
rect 28215 35680 28227 35683
rect 28902 35680 28908 35692
rect 28215 35652 28908 35680
rect 28215 35649 28227 35652
rect 28169 35643 28227 35649
rect 28902 35640 28908 35652
rect 28960 35640 28966 35692
rect 23750 35612 23756 35624
rect 22204 35584 23756 35612
rect 23750 35572 23756 35584
rect 23808 35572 23814 35624
rect 24026 35612 24032 35624
rect 23987 35584 24032 35612
rect 24026 35572 24032 35584
rect 24084 35572 24090 35624
rect 27706 35612 27712 35624
rect 27667 35584 27712 35612
rect 27706 35572 27712 35584
rect 27764 35572 27770 35624
rect 27801 35615 27859 35621
rect 27801 35581 27813 35615
rect 27847 35581 27859 35615
rect 28994 35612 29000 35624
rect 27801 35575 27859 35581
rect 28184 35584 29000 35612
rect 14921 35547 14979 35553
rect 14921 35544 14933 35547
rect 13596 35516 14933 35544
rect 13596 35504 13602 35516
rect 14921 35513 14933 35516
rect 14967 35513 14979 35547
rect 14921 35507 14979 35513
rect 20533 35547 20591 35553
rect 20533 35513 20545 35547
rect 20579 35513 20591 35547
rect 27816 35544 27844 35575
rect 28184 35544 28212 35584
rect 28994 35572 29000 35584
rect 29052 35612 29058 35624
rect 29730 35612 29736 35624
rect 29052 35584 29736 35612
rect 29052 35572 29058 35584
rect 29730 35572 29736 35584
rect 29788 35572 29794 35624
rect 30484 35612 30512 35720
rect 31202 35708 31208 35720
rect 31260 35708 31266 35760
rect 31573 35751 31631 35757
rect 31573 35717 31585 35751
rect 31619 35748 31631 35751
rect 32585 35751 32643 35757
rect 32585 35748 32597 35751
rect 31619 35720 32597 35748
rect 31619 35717 31631 35720
rect 31573 35711 31631 35717
rect 32585 35717 32597 35720
rect 32631 35717 32643 35751
rect 32585 35711 32643 35717
rect 30834 35680 30840 35692
rect 30747 35652 30840 35680
rect 30834 35640 30840 35652
rect 30892 35680 30898 35692
rect 31481 35683 31539 35689
rect 31481 35680 31493 35683
rect 30892 35652 31493 35680
rect 30892 35640 30898 35652
rect 31481 35649 31493 35652
rect 31527 35649 31539 35683
rect 31481 35643 31539 35649
rect 31665 35683 31723 35689
rect 31665 35649 31677 35683
rect 31711 35649 31723 35683
rect 32306 35680 32312 35692
rect 32267 35652 32312 35680
rect 31665 35643 31723 35649
rect 30116 35584 30512 35612
rect 27816 35516 28212 35544
rect 20533 35507 20591 35513
rect 28626 35504 28632 35556
rect 28684 35544 28690 35556
rect 29089 35547 29147 35553
rect 29089 35544 29101 35547
rect 28684 35516 29101 35544
rect 28684 35504 28690 35516
rect 29089 35513 29101 35516
rect 29135 35513 29147 35547
rect 30116 35544 30144 35584
rect 30558 35572 30564 35624
rect 30616 35612 30622 35624
rect 30653 35615 30711 35621
rect 30653 35612 30665 35615
rect 30616 35584 30665 35612
rect 30616 35572 30622 35584
rect 30653 35581 30665 35584
rect 30699 35581 30711 35615
rect 30653 35575 30711 35581
rect 29089 35507 29147 35513
rect 30024 35516 30144 35544
rect 30193 35547 30251 35553
rect 14458 35476 14464 35488
rect 9640 35448 12112 35476
rect 14419 35448 14464 35476
rect 9640 35436 9646 35448
rect 14458 35436 14464 35448
rect 14516 35436 14522 35488
rect 16114 35476 16120 35488
rect 16075 35448 16120 35476
rect 16114 35436 16120 35448
rect 16172 35436 16178 35488
rect 16390 35436 16396 35488
rect 16448 35476 16454 35488
rect 17497 35479 17555 35485
rect 17497 35476 17509 35479
rect 16448 35448 17509 35476
rect 16448 35436 16454 35448
rect 17497 35445 17509 35448
rect 17543 35445 17555 35479
rect 17497 35439 17555 35445
rect 20898 35436 20904 35488
rect 20956 35476 20962 35488
rect 20993 35479 21051 35485
rect 20993 35476 21005 35479
rect 20956 35448 21005 35476
rect 20956 35436 20962 35448
rect 20993 35445 21005 35448
rect 21039 35445 21051 35479
rect 20993 35439 21051 35445
rect 22002 35436 22008 35488
rect 22060 35476 22066 35488
rect 22097 35479 22155 35485
rect 22097 35476 22109 35479
rect 22060 35448 22109 35476
rect 22060 35436 22066 35448
rect 22097 35445 22109 35448
rect 22143 35445 22155 35479
rect 22738 35476 22744 35488
rect 22699 35448 22744 35476
rect 22097 35439 22155 35445
rect 22738 35436 22744 35448
rect 22796 35436 22802 35488
rect 28350 35476 28356 35488
rect 28311 35448 28356 35476
rect 28350 35436 28356 35448
rect 28408 35436 28414 35488
rect 29273 35479 29331 35485
rect 29273 35445 29285 35479
rect 29319 35476 29331 35479
rect 29362 35476 29368 35488
rect 29319 35448 29368 35476
rect 29319 35445 29331 35448
rect 29273 35439 29331 35445
rect 29362 35436 29368 35448
rect 29420 35436 29426 35488
rect 30024 35485 30052 35516
rect 30193 35513 30205 35547
rect 30239 35544 30251 35547
rect 30852 35544 30880 35640
rect 30926 35572 30932 35624
rect 30984 35612 30990 35624
rect 31680 35612 31708 35643
rect 32306 35640 32312 35652
rect 32364 35640 32370 35692
rect 33686 35640 33692 35692
rect 33744 35640 33750 35692
rect 30984 35584 31708 35612
rect 30984 35572 30990 35584
rect 30239 35516 30880 35544
rect 30239 35513 30251 35516
rect 30193 35507 30251 35513
rect 30009 35479 30067 35485
rect 30009 35445 30021 35479
rect 30055 35445 30067 35479
rect 30009 35439 30067 35445
rect 30098 35436 30104 35488
rect 30156 35476 30162 35488
rect 31021 35479 31079 35485
rect 31021 35476 31033 35479
rect 30156 35448 31033 35476
rect 30156 35436 30162 35448
rect 31021 35445 31033 35448
rect 31067 35476 31079 35479
rect 31478 35476 31484 35488
rect 31067 35448 31484 35476
rect 31067 35445 31079 35448
rect 31021 35439 31079 35445
rect 31478 35436 31484 35448
rect 31536 35436 31542 35488
rect 1104 35386 37628 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 37628 35386
rect 1104 35312 37628 35334
rect 6730 35232 6736 35284
rect 6788 35272 6794 35284
rect 6898 35275 6956 35281
rect 6898 35272 6910 35275
rect 6788 35244 6910 35272
rect 6788 35232 6794 35244
rect 6898 35241 6910 35244
rect 6944 35241 6956 35275
rect 6898 35235 6956 35241
rect 8110 35232 8116 35284
rect 8168 35272 8174 35284
rect 8389 35275 8447 35281
rect 8389 35272 8401 35275
rect 8168 35244 8401 35272
rect 8168 35232 8174 35244
rect 8389 35241 8401 35244
rect 8435 35241 8447 35275
rect 10318 35272 10324 35284
rect 10279 35244 10324 35272
rect 8389 35235 8447 35241
rect 6641 35139 6699 35145
rect 6641 35105 6653 35139
rect 6687 35136 6699 35139
rect 8202 35136 8208 35148
rect 6687 35108 8208 35136
rect 6687 35105 6699 35108
rect 6641 35099 6699 35105
rect 8202 35096 8208 35108
rect 8260 35096 8266 35148
rect 8404 35136 8432 35235
rect 10318 35232 10324 35244
rect 10376 35232 10382 35284
rect 17954 35232 17960 35284
rect 18012 35272 18018 35284
rect 18233 35275 18291 35281
rect 18233 35272 18245 35275
rect 18012 35244 18245 35272
rect 18012 35232 18018 35244
rect 18233 35241 18245 35244
rect 18279 35241 18291 35275
rect 21358 35272 21364 35284
rect 18233 35235 18291 35241
rect 20548 35244 21364 35272
rect 12158 35204 12164 35216
rect 9784 35176 12164 35204
rect 9784 35145 9812 35176
rect 10336 35148 10364 35176
rect 12158 35164 12164 35176
rect 12216 35164 12222 35216
rect 9585 35139 9643 35145
rect 9585 35136 9597 35139
rect 8404 35108 9597 35136
rect 9585 35105 9597 35108
rect 9631 35105 9643 35139
rect 9585 35099 9643 35105
rect 9769 35139 9827 35145
rect 9769 35105 9781 35139
rect 9815 35105 9827 35139
rect 9769 35099 9827 35105
rect 1765 35071 1823 35077
rect 1765 35037 1777 35071
rect 1811 35068 1823 35071
rect 2038 35068 2044 35080
rect 1811 35040 2044 35068
rect 1811 35037 1823 35040
rect 1765 35031 1823 35037
rect 2038 35028 2044 35040
rect 2096 35028 2102 35080
rect 9600 35068 9628 35099
rect 10318 35096 10324 35148
rect 10376 35096 10382 35148
rect 10594 35096 10600 35148
rect 10652 35136 10658 35148
rect 10962 35136 10968 35148
rect 10652 35108 10968 35136
rect 10652 35096 10658 35108
rect 10962 35096 10968 35108
rect 11020 35096 11026 35148
rect 13814 35096 13820 35148
rect 13872 35136 13878 35148
rect 14277 35139 14335 35145
rect 14277 35136 14289 35139
rect 13872 35108 14289 35136
rect 13872 35096 13878 35108
rect 14277 35105 14289 35108
rect 14323 35136 14335 35139
rect 14550 35136 14556 35148
rect 14323 35108 14556 35136
rect 14323 35105 14335 35108
rect 14277 35099 14335 35105
rect 14550 35096 14556 35108
rect 14608 35096 14614 35148
rect 16485 35139 16543 35145
rect 16485 35105 16497 35139
rect 16531 35136 16543 35139
rect 16758 35136 16764 35148
rect 16531 35108 16764 35136
rect 16531 35105 16543 35108
rect 16485 35099 16543 35105
rect 16758 35096 16764 35108
rect 16816 35136 16822 35148
rect 17310 35136 17316 35148
rect 16816 35108 17316 35136
rect 16816 35096 16822 35108
rect 17310 35096 17316 35108
rect 17368 35096 17374 35148
rect 19886 35136 19892 35148
rect 19847 35108 19892 35136
rect 19886 35096 19892 35108
rect 19944 35096 19950 35148
rect 19978 35096 19984 35148
rect 20036 35136 20042 35148
rect 20346 35136 20352 35148
rect 20036 35108 20352 35136
rect 20036 35096 20042 35108
rect 20346 35096 20352 35108
rect 20404 35096 20410 35148
rect 10781 35071 10839 35077
rect 10781 35068 10793 35071
rect 9600 35040 10793 35068
rect 10781 35037 10793 35040
rect 10827 35037 10839 35071
rect 10781 35031 10839 35037
rect 11609 35071 11667 35077
rect 11609 35037 11621 35071
rect 11655 35068 11667 35071
rect 12158 35068 12164 35080
rect 11655 35040 12164 35068
rect 11655 35037 11667 35040
rect 11609 35031 11667 35037
rect 12158 35028 12164 35040
rect 12216 35028 12222 35080
rect 12253 35071 12311 35077
rect 12253 35037 12265 35071
rect 12299 35037 12311 35071
rect 12253 35031 12311 35037
rect 7374 34960 7380 35012
rect 7432 34960 7438 35012
rect 11238 34960 11244 35012
rect 11296 35000 11302 35012
rect 12268 35000 12296 35031
rect 12434 35028 12440 35080
rect 12492 35068 12498 35080
rect 12618 35068 12624 35080
rect 12492 35040 12624 35068
rect 12492 35028 12498 35040
rect 12618 35028 12624 35040
rect 12676 35068 12682 35080
rect 12897 35071 12955 35077
rect 12897 35068 12909 35071
rect 12676 35040 12909 35068
rect 12676 35028 12682 35040
rect 12897 35037 12909 35040
rect 12943 35037 12955 35071
rect 13538 35068 13544 35080
rect 13499 35040 13544 35068
rect 12897 35031 12955 35037
rect 13538 35028 13544 35040
rect 13596 35028 13602 35080
rect 18877 35071 18935 35077
rect 18877 35037 18889 35071
rect 18923 35068 18935 35071
rect 19242 35068 19248 35080
rect 18923 35040 19248 35068
rect 18923 35037 18935 35040
rect 18877 35031 18935 35037
rect 19242 35028 19248 35040
rect 19300 35068 19306 35080
rect 20548 35068 20576 35244
rect 21358 35232 21364 35244
rect 21416 35232 21422 35284
rect 22370 35272 22376 35284
rect 22331 35244 22376 35272
rect 22370 35232 22376 35244
rect 22428 35232 22434 35284
rect 23290 35272 23296 35284
rect 23251 35244 23296 35272
rect 23290 35232 23296 35244
rect 23348 35232 23354 35284
rect 27249 35275 27307 35281
rect 27249 35241 27261 35275
rect 27295 35272 27307 35275
rect 27614 35272 27620 35284
rect 27295 35244 27620 35272
rect 27295 35241 27307 35244
rect 27249 35235 27307 35241
rect 27614 35232 27620 35244
rect 27672 35232 27678 35284
rect 28166 35272 28172 35284
rect 28127 35244 28172 35272
rect 28166 35232 28172 35244
rect 28224 35232 28230 35284
rect 28353 35275 28411 35281
rect 28353 35241 28365 35275
rect 28399 35272 28411 35275
rect 28534 35272 28540 35284
rect 28399 35244 28540 35272
rect 28399 35241 28411 35244
rect 28353 35235 28411 35241
rect 28534 35232 28540 35244
rect 28592 35232 28598 35284
rect 28629 35275 28687 35281
rect 28629 35241 28641 35275
rect 28675 35272 28687 35275
rect 28810 35272 28816 35284
rect 28675 35244 28816 35272
rect 28675 35241 28687 35244
rect 28629 35235 28687 35241
rect 28810 35232 28816 35244
rect 28868 35232 28874 35284
rect 29914 35272 29920 35284
rect 29875 35244 29920 35272
rect 29914 35232 29920 35244
rect 29972 35232 29978 35284
rect 33042 35232 33048 35284
rect 33100 35272 33106 35284
rect 33505 35275 33563 35281
rect 33505 35272 33517 35275
rect 33100 35244 33517 35272
rect 33100 35232 33106 35244
rect 33505 35241 33517 35244
rect 33551 35241 33563 35275
rect 33505 35235 33563 35241
rect 22186 35164 22192 35216
rect 22244 35204 22250 35216
rect 26970 35204 26976 35216
rect 22244 35176 26976 35204
rect 22244 35164 22250 35176
rect 26970 35164 26976 35176
rect 27028 35164 27034 35216
rect 20625 35139 20683 35145
rect 20625 35105 20637 35139
rect 20671 35136 20683 35139
rect 22094 35136 22100 35148
rect 20671 35108 22100 35136
rect 20671 35105 20683 35108
rect 20625 35099 20683 35105
rect 22094 35096 22100 35108
rect 22152 35096 22158 35148
rect 23382 35096 23388 35148
rect 23440 35136 23446 35148
rect 23566 35136 23572 35148
rect 23440 35108 23572 35136
rect 23440 35096 23446 35108
rect 23566 35096 23572 35108
rect 23624 35136 23630 35148
rect 23845 35139 23903 35145
rect 23845 35136 23857 35139
rect 23624 35108 23857 35136
rect 23624 35096 23630 35108
rect 23845 35105 23857 35108
rect 23891 35105 23903 35139
rect 23845 35099 23903 35105
rect 24765 35139 24823 35145
rect 24765 35105 24777 35139
rect 24811 35136 24823 35139
rect 25038 35136 25044 35148
rect 24811 35108 25044 35136
rect 24811 35105 24823 35108
rect 24765 35099 24823 35105
rect 25038 35096 25044 35108
rect 25096 35096 25102 35148
rect 26050 35096 26056 35148
rect 26108 35136 26114 35148
rect 26329 35139 26387 35145
rect 26329 35136 26341 35139
rect 26108 35108 26341 35136
rect 26108 35096 26114 35108
rect 26329 35105 26341 35108
rect 26375 35105 26387 35139
rect 26329 35099 26387 35105
rect 19300 35040 20576 35068
rect 19300 35028 19306 35040
rect 22002 35028 22008 35080
rect 22060 35028 22066 35080
rect 24949 35071 25007 35077
rect 24949 35037 24961 35071
rect 24995 35068 25007 35071
rect 26237 35071 26295 35077
rect 26237 35068 26249 35071
rect 24995 35040 26249 35068
rect 24995 35037 25007 35040
rect 24949 35031 25007 35037
rect 26237 35037 26249 35040
rect 26283 35068 26295 35071
rect 26694 35068 26700 35080
rect 26283 35040 26700 35068
rect 26283 35037 26295 35040
rect 26237 35031 26295 35037
rect 26694 35028 26700 35040
rect 26752 35028 26758 35080
rect 26988 35077 27016 35164
rect 27246 35096 27252 35148
rect 27304 35136 27310 35148
rect 28258 35136 28264 35148
rect 27304 35108 28120 35136
rect 28219 35108 28264 35136
rect 27304 35096 27310 35108
rect 26973 35071 27031 35077
rect 26973 35037 26985 35071
rect 27019 35037 27031 35071
rect 27890 35068 27896 35080
rect 27851 35040 27896 35068
rect 26973 35031 27031 35037
rect 27890 35028 27896 35040
rect 27948 35028 27954 35080
rect 28092 35077 28120 35108
rect 28258 35096 28264 35108
rect 28316 35096 28322 35148
rect 32306 35096 32312 35148
rect 32364 35136 32370 35148
rect 32953 35139 33011 35145
rect 32953 35136 32965 35139
rect 32364 35108 32965 35136
rect 32364 35096 32370 35108
rect 32953 35105 32965 35108
rect 32999 35105 33011 35139
rect 32953 35099 33011 35105
rect 28077 35071 28135 35077
rect 28077 35037 28089 35071
rect 28123 35037 28135 35071
rect 28077 35031 28135 35037
rect 13446 35000 13452 35012
rect 11296 34972 13452 35000
rect 11296 34960 11302 34972
rect 13446 34960 13452 34972
rect 13504 34960 13510 35012
rect 14553 35003 14611 35009
rect 14553 35000 14565 35003
rect 13740 34972 14565 35000
rect 1578 34932 1584 34944
rect 1539 34904 1584 34932
rect 1578 34892 1584 34904
rect 1636 34892 1642 34944
rect 8846 34892 8852 34944
rect 8904 34932 8910 34944
rect 9125 34935 9183 34941
rect 9125 34932 9137 34935
rect 8904 34904 9137 34932
rect 8904 34892 8910 34904
rect 9125 34901 9137 34904
rect 9171 34901 9183 34935
rect 9490 34932 9496 34944
rect 9451 34904 9496 34932
rect 9125 34895 9183 34901
rect 9490 34892 9496 34904
rect 9548 34892 9554 34944
rect 10594 34892 10600 34944
rect 10652 34932 10658 34944
rect 10689 34935 10747 34941
rect 10689 34932 10701 34935
rect 10652 34904 10701 34932
rect 10652 34892 10658 34904
rect 10689 34901 10701 34904
rect 10735 34901 10747 34935
rect 11790 34932 11796 34944
rect 11751 34904 11796 34932
rect 10689 34895 10747 34901
rect 11790 34892 11796 34904
rect 11848 34892 11854 34944
rect 12342 34932 12348 34944
rect 12303 34904 12348 34932
rect 12342 34892 12348 34904
rect 12400 34892 12406 34944
rect 12986 34932 12992 34944
rect 12947 34904 12992 34932
rect 12986 34892 12992 34904
rect 13044 34892 13050 34944
rect 13740 34941 13768 34972
rect 14553 34969 14565 34972
rect 14599 34969 14611 35003
rect 14553 34963 14611 34969
rect 15562 34960 15568 35012
rect 15620 34960 15626 35012
rect 16298 34960 16304 35012
rect 16356 35000 16362 35012
rect 16761 35003 16819 35009
rect 16761 35000 16773 35003
rect 16356 34972 16773 35000
rect 16356 34960 16362 34972
rect 16761 34969 16773 34972
rect 16807 34969 16819 35003
rect 18785 35003 18843 35009
rect 18785 35000 18797 35003
rect 17986 34972 18797 35000
rect 16761 34963 16819 34969
rect 18785 34969 18797 34972
rect 18831 34969 18843 35003
rect 18785 34963 18843 34969
rect 19518 34960 19524 35012
rect 19576 35000 19582 35012
rect 20898 35000 20904 35012
rect 19576 34972 20760 35000
rect 20859 34972 20904 35000
rect 19576 34960 19582 34972
rect 13725 34935 13783 34941
rect 13725 34901 13737 34935
rect 13771 34901 13783 34935
rect 13725 34895 13783 34901
rect 15930 34892 15936 34944
rect 15988 34932 15994 34944
rect 16025 34935 16083 34941
rect 16025 34932 16037 34935
rect 15988 34904 16037 34932
rect 15988 34892 15994 34904
rect 16025 34901 16037 34904
rect 16071 34901 16083 34935
rect 16025 34895 16083 34901
rect 19334 34892 19340 34944
rect 19392 34932 19398 34944
rect 19429 34935 19487 34941
rect 19429 34932 19441 34935
rect 19392 34904 19441 34932
rect 19392 34892 19398 34904
rect 19429 34901 19441 34904
rect 19475 34901 19487 34935
rect 19794 34932 19800 34944
rect 19755 34904 19800 34932
rect 19429 34895 19487 34901
rect 19794 34892 19800 34904
rect 19852 34892 19858 34944
rect 20732 34932 20760 34972
rect 20898 34960 20904 34972
rect 20956 34960 20962 35012
rect 23661 35003 23719 35009
rect 23661 34969 23673 35003
rect 23707 35000 23719 35003
rect 26142 35000 26148 35012
rect 23707 34972 25820 35000
rect 26103 34972 26148 35000
rect 23707 34969 23719 34972
rect 23661 34963 23719 34969
rect 23382 34932 23388 34944
rect 20732 34904 23388 34932
rect 23382 34892 23388 34904
rect 23440 34892 23446 34944
rect 23753 34935 23811 34941
rect 23753 34901 23765 34935
rect 23799 34932 23811 34935
rect 23934 34932 23940 34944
rect 23799 34904 23940 34932
rect 23799 34901 23811 34904
rect 23753 34895 23811 34901
rect 23934 34892 23940 34904
rect 23992 34932 23998 34944
rect 24857 34935 24915 34941
rect 24857 34932 24869 34935
rect 23992 34904 24869 34932
rect 23992 34892 23998 34904
rect 24857 34901 24869 34904
rect 24903 34901 24915 34935
rect 24857 34895 24915 34901
rect 25317 34935 25375 34941
rect 25317 34901 25329 34935
rect 25363 34932 25375 34935
rect 25682 34932 25688 34944
rect 25363 34904 25688 34932
rect 25363 34901 25375 34904
rect 25317 34895 25375 34901
rect 25682 34892 25688 34904
rect 25740 34892 25746 34944
rect 25792 34941 25820 34972
rect 26142 34960 26148 34972
rect 26200 34960 26206 35012
rect 28276 35000 28304 35096
rect 28442 35028 28448 35080
rect 28500 35068 28506 35080
rect 30193 35071 30251 35077
rect 30193 35068 30205 35071
rect 28500 35040 30205 35068
rect 28500 35028 28506 35040
rect 30193 35037 30205 35040
rect 30239 35037 30251 35071
rect 30193 35031 30251 35037
rect 33502 35028 33508 35080
rect 33560 35068 33566 35080
rect 33597 35071 33655 35077
rect 33597 35068 33609 35071
rect 33560 35040 33609 35068
rect 33560 35028 33566 35040
rect 33597 35037 33609 35040
rect 33643 35037 33655 35071
rect 36906 35068 36912 35080
rect 36867 35040 36912 35068
rect 33597 35031 33655 35037
rect 36906 35028 36912 35040
rect 36964 35028 36970 35080
rect 28534 35000 28540 35012
rect 28276 34972 28540 35000
rect 28534 34960 28540 34972
rect 28592 34960 28598 35012
rect 32674 35000 32680 35012
rect 32246 34972 32536 35000
rect 32635 34972 32680 35000
rect 25777 34935 25835 34941
rect 25777 34901 25789 34935
rect 25823 34901 25835 34935
rect 25777 34895 25835 34901
rect 27433 34935 27491 34941
rect 27433 34901 27445 34935
rect 27479 34932 27491 34935
rect 28258 34932 28264 34944
rect 27479 34904 28264 34932
rect 27479 34901 27491 34904
rect 27433 34895 27491 34901
rect 28258 34892 28264 34904
rect 28316 34892 28322 34944
rect 28442 34892 28448 34944
rect 28500 34932 28506 34944
rect 29733 34935 29791 34941
rect 29733 34932 29745 34935
rect 28500 34904 29745 34932
rect 28500 34892 28506 34904
rect 29733 34901 29745 34904
rect 29779 34901 29791 34935
rect 29733 34895 29791 34901
rect 30558 34892 30564 34944
rect 30616 34932 30622 34944
rect 31205 34935 31263 34941
rect 31205 34932 31217 34935
rect 30616 34904 31217 34932
rect 30616 34892 30622 34904
rect 31205 34901 31217 34904
rect 31251 34901 31263 34935
rect 32508 34932 32536 34972
rect 32674 34960 32680 34972
rect 32732 34960 32738 35012
rect 33134 34932 33140 34944
rect 32508 34904 33140 34932
rect 31205 34895 31263 34901
rect 33134 34892 33140 34904
rect 33192 34892 33198 34944
rect 37090 34932 37096 34944
rect 37051 34904 37096 34932
rect 37090 34892 37096 34904
rect 37148 34892 37154 34944
rect 1104 34842 37628 34864
rect 1104 34790 4874 34842
rect 4926 34790 4938 34842
rect 4990 34790 5002 34842
rect 5054 34790 5066 34842
rect 5118 34790 5130 34842
rect 5182 34790 35594 34842
rect 35646 34790 35658 34842
rect 35710 34790 35722 34842
rect 35774 34790 35786 34842
rect 35838 34790 35850 34842
rect 35902 34790 37628 34842
rect 1104 34768 37628 34790
rect 7190 34688 7196 34740
rect 7248 34728 7254 34740
rect 8481 34731 8539 34737
rect 8481 34728 8493 34731
rect 7248 34700 8493 34728
rect 7248 34688 7254 34700
rect 8481 34697 8493 34700
rect 8527 34697 8539 34731
rect 8846 34728 8852 34740
rect 8807 34700 8852 34728
rect 8481 34691 8539 34697
rect 8846 34688 8852 34700
rect 8904 34688 8910 34740
rect 8941 34731 8999 34737
rect 8941 34697 8953 34731
rect 8987 34728 8999 34731
rect 9582 34728 9588 34740
rect 8987 34700 9588 34728
rect 8987 34697 8999 34700
rect 8941 34691 8999 34697
rect 9582 34688 9588 34700
rect 9640 34688 9646 34740
rect 11701 34731 11759 34737
rect 11701 34697 11713 34731
rect 11747 34697 11759 34731
rect 11701 34691 11759 34697
rect 12989 34731 13047 34737
rect 12989 34697 13001 34731
rect 13035 34728 13047 34731
rect 13170 34728 13176 34740
rect 13035 34700 13176 34728
rect 13035 34697 13047 34700
rect 12989 34691 13047 34697
rect 11716 34660 11744 34691
rect 13170 34688 13176 34700
rect 13228 34688 13234 34740
rect 13446 34688 13452 34740
rect 13504 34728 13510 34740
rect 15562 34728 15568 34740
rect 13504 34700 14872 34728
rect 15523 34700 15568 34728
rect 13504 34688 13510 34700
rect 10336 34632 11744 34660
rect 10336 34601 10364 34632
rect 12342 34620 12348 34672
rect 12400 34660 12406 34672
rect 12400 34632 13294 34660
rect 12400 34620 12406 34632
rect 14550 34620 14556 34672
rect 14608 34660 14614 34672
rect 14844 34660 14872 34700
rect 15562 34688 15568 34700
rect 15620 34688 15626 34740
rect 16298 34728 16304 34740
rect 16259 34700 16304 34728
rect 16298 34688 16304 34700
rect 16356 34688 16362 34740
rect 17862 34688 17868 34740
rect 17920 34728 17926 34740
rect 18049 34731 18107 34737
rect 18049 34728 18061 34731
rect 17920 34700 18061 34728
rect 17920 34688 17926 34700
rect 18049 34697 18061 34700
rect 18095 34697 18107 34731
rect 18049 34691 18107 34697
rect 18509 34731 18567 34737
rect 18509 34697 18521 34731
rect 18555 34728 18567 34731
rect 18598 34728 18604 34740
rect 18555 34700 18604 34728
rect 18555 34697 18567 34700
rect 18509 34691 18567 34697
rect 18598 34688 18604 34700
rect 18656 34688 18662 34740
rect 23934 34728 23940 34740
rect 23895 34700 23940 34728
rect 23934 34688 23940 34700
rect 23992 34728 23998 34740
rect 24765 34731 24823 34737
rect 24765 34728 24777 34731
rect 23992 34700 24777 34728
rect 23992 34688 23998 34700
rect 24765 34697 24777 34700
rect 24811 34697 24823 34731
rect 24765 34691 24823 34697
rect 24857 34731 24915 34737
rect 24857 34697 24869 34731
rect 24903 34728 24915 34731
rect 24946 34728 24952 34740
rect 24903 34700 24952 34728
rect 24903 34697 24915 34700
rect 24857 34691 24915 34697
rect 24946 34688 24952 34700
rect 25004 34688 25010 34740
rect 25685 34731 25743 34737
rect 25685 34697 25697 34731
rect 25731 34697 25743 34731
rect 28258 34728 28264 34740
rect 28219 34700 28264 34728
rect 25685 34691 25743 34697
rect 22465 34663 22523 34669
rect 14608 34632 14780 34660
rect 14844 34632 17448 34660
rect 14608 34620 14614 34632
rect 10321 34595 10379 34601
rect 10321 34561 10333 34595
rect 10367 34561 10379 34595
rect 10321 34555 10379 34561
rect 10965 34595 11023 34601
rect 10965 34561 10977 34595
rect 11011 34592 11023 34595
rect 11238 34592 11244 34604
rect 11011 34564 11244 34592
rect 11011 34561 11023 34564
rect 10965 34555 11023 34561
rect 11238 34552 11244 34564
rect 11296 34552 11302 34604
rect 12066 34592 12072 34604
rect 12027 34564 12072 34592
rect 12066 34552 12072 34564
rect 12124 34552 12130 34604
rect 14752 34601 14780 34632
rect 15672 34601 15700 34632
rect 14737 34595 14795 34601
rect 14737 34561 14749 34595
rect 14783 34561 14795 34595
rect 14737 34555 14795 34561
rect 15657 34595 15715 34601
rect 15657 34561 15669 34595
rect 15703 34561 15715 34595
rect 15657 34555 15715 34561
rect 16117 34595 16175 34601
rect 16117 34561 16129 34595
rect 16163 34592 16175 34595
rect 16390 34592 16396 34604
rect 16163 34564 16396 34592
rect 16163 34561 16175 34564
rect 16117 34555 16175 34561
rect 16390 34552 16396 34564
rect 16448 34552 16454 34604
rect 17420 34601 17448 34632
rect 22465 34629 22477 34663
rect 22511 34660 22523 34663
rect 22738 34660 22744 34672
rect 22511 34632 22744 34660
rect 22511 34629 22523 34632
rect 22465 34623 22523 34629
rect 22738 34620 22744 34632
rect 22796 34620 22802 34672
rect 25700 34660 25728 34691
rect 28258 34688 28264 34700
rect 28316 34688 28322 34740
rect 28626 34728 28632 34740
rect 28587 34700 28632 34728
rect 28626 34688 28632 34700
rect 28684 34688 28690 34740
rect 29914 34688 29920 34740
rect 29972 34688 29978 34740
rect 30926 34737 30932 34740
rect 30922 34728 30932 34737
rect 30887 34700 30932 34728
rect 30922 34691 30932 34700
rect 30926 34688 30932 34691
rect 30984 34688 30990 34740
rect 31573 34731 31631 34737
rect 31573 34697 31585 34731
rect 31619 34728 31631 34731
rect 32674 34728 32680 34740
rect 31619 34700 32680 34728
rect 31619 34697 31631 34700
rect 31573 34691 31631 34697
rect 32674 34688 32680 34700
rect 32732 34688 32738 34740
rect 23690 34632 25728 34660
rect 28169 34663 28227 34669
rect 28169 34629 28181 34663
rect 28215 34660 28227 34663
rect 28442 34660 28448 34672
rect 28215 34632 28448 34660
rect 28215 34629 28227 34632
rect 28169 34623 28227 34629
rect 28442 34620 28448 34632
rect 28500 34620 28506 34672
rect 29932 34660 29960 34688
rect 31021 34663 31079 34669
rect 31021 34660 31033 34663
rect 29288 34632 31033 34660
rect 17405 34595 17463 34601
rect 17405 34561 17417 34595
rect 17451 34592 17463 34595
rect 18046 34592 18052 34604
rect 17451 34564 18052 34592
rect 17451 34561 17463 34564
rect 17405 34555 17463 34561
rect 18046 34552 18052 34564
rect 18104 34552 18110 34604
rect 18414 34592 18420 34604
rect 18375 34564 18420 34592
rect 18414 34552 18420 34564
rect 18472 34552 18478 34604
rect 19426 34592 19432 34604
rect 19387 34564 19432 34592
rect 19426 34552 19432 34564
rect 19484 34552 19490 34604
rect 20806 34552 20812 34604
rect 20864 34552 20870 34604
rect 23750 34552 23756 34604
rect 23808 34592 23814 34604
rect 25593 34595 25651 34601
rect 25593 34592 25605 34595
rect 23808 34564 25605 34592
rect 23808 34552 23814 34564
rect 25593 34561 25605 34564
rect 25639 34561 25651 34595
rect 25593 34555 25651 34561
rect 25682 34552 25688 34604
rect 25740 34592 25746 34604
rect 26421 34595 26479 34601
rect 26421 34592 26433 34595
rect 25740 34564 26433 34592
rect 25740 34552 25746 34564
rect 26421 34561 26433 34564
rect 26467 34561 26479 34595
rect 26421 34555 26479 34561
rect 27246 34552 27252 34604
rect 27304 34592 27310 34604
rect 27893 34595 27951 34601
rect 27893 34592 27905 34595
rect 27304 34564 27905 34592
rect 27304 34552 27310 34564
rect 27893 34561 27905 34564
rect 27939 34561 27951 34595
rect 27893 34555 27951 34561
rect 28353 34595 28411 34601
rect 28353 34561 28365 34595
rect 28399 34592 28411 34595
rect 28994 34592 29000 34604
rect 28399 34564 29000 34592
rect 28399 34561 28411 34564
rect 28353 34555 28411 34561
rect 28994 34552 29000 34564
rect 29052 34552 29058 34604
rect 29288 34601 29316 34632
rect 31021 34629 31033 34632
rect 31067 34629 31079 34663
rect 31021 34623 31079 34629
rect 31110 34620 31116 34672
rect 31168 34660 31174 34672
rect 32309 34663 32367 34669
rect 32309 34660 32321 34663
rect 31168 34632 32321 34660
rect 31168 34620 31174 34632
rect 32309 34629 32321 34632
rect 32355 34629 32367 34663
rect 32309 34623 32367 34629
rect 29273 34595 29331 34601
rect 29273 34561 29285 34595
rect 29319 34561 29331 34595
rect 29914 34592 29920 34604
rect 29875 34564 29920 34592
rect 29273 34555 29331 34561
rect 29914 34552 29920 34564
rect 29972 34552 29978 34604
rect 30745 34595 30803 34601
rect 30745 34592 30757 34595
rect 30392 34564 30757 34592
rect 30392 34536 30420 34564
rect 30745 34561 30757 34564
rect 30791 34561 30803 34595
rect 30745 34555 30803 34561
rect 30837 34595 30895 34601
rect 30837 34561 30849 34595
rect 30883 34592 30895 34595
rect 31202 34592 31208 34604
rect 30883 34564 31208 34592
rect 30883 34561 30895 34564
rect 30837 34555 30895 34561
rect 9125 34527 9183 34533
rect 9125 34493 9137 34527
rect 9171 34493 9183 34527
rect 9125 34487 9183 34493
rect 9140 34456 9168 34487
rect 10686 34484 10692 34536
rect 10744 34484 10750 34536
rect 11057 34527 11115 34533
rect 11057 34493 11069 34527
rect 11103 34524 11115 34527
rect 11146 34524 11152 34536
rect 11103 34496 11152 34524
rect 11103 34493 11115 34496
rect 11057 34487 11115 34493
rect 11146 34484 11152 34496
rect 11204 34484 11210 34536
rect 11974 34484 11980 34536
rect 12032 34524 12038 34536
rect 12161 34527 12219 34533
rect 12161 34524 12173 34527
rect 12032 34496 12173 34524
rect 12032 34484 12038 34496
rect 12161 34493 12173 34496
rect 12207 34493 12219 34527
rect 12161 34487 12219 34493
rect 12345 34527 12403 34533
rect 12345 34493 12357 34527
rect 12391 34524 12403 34527
rect 13906 34524 13912 34536
rect 12391 34496 13912 34524
rect 12391 34493 12403 34496
rect 12345 34487 12403 34493
rect 9674 34456 9680 34468
rect 9140 34428 9680 34456
rect 9674 34416 9680 34428
rect 9732 34456 9738 34468
rect 10704 34456 10732 34484
rect 10870 34456 10876 34468
rect 9732 34428 10876 34456
rect 9732 34416 9738 34428
rect 10870 34416 10876 34428
rect 10928 34456 10934 34468
rect 12360 34456 12388 34487
rect 13906 34484 13912 34496
rect 13964 34484 13970 34536
rect 18601 34527 18659 34533
rect 18601 34493 18613 34527
rect 18647 34493 18659 34527
rect 18601 34487 18659 34493
rect 10928 34428 12388 34456
rect 10928 34416 10934 34428
rect 16022 34416 16028 34468
rect 16080 34456 16086 34468
rect 18616 34456 18644 34487
rect 19794 34484 19800 34536
rect 19852 34524 19858 34536
rect 21177 34527 21235 34533
rect 21177 34524 21189 34527
rect 19852 34496 21189 34524
rect 19852 34484 19858 34496
rect 21177 34493 21189 34496
rect 21223 34524 21235 34527
rect 21223 34496 22048 34524
rect 21223 34493 21235 34496
rect 21177 34487 21235 34493
rect 16080 34428 18644 34456
rect 22020 34456 22048 34496
rect 22094 34484 22100 34536
rect 22152 34524 22158 34536
rect 22189 34527 22247 34533
rect 22189 34524 22201 34527
rect 22152 34496 22201 34524
rect 22152 34484 22158 34496
rect 22189 34493 22201 34496
rect 22235 34524 22247 34527
rect 22235 34496 23520 34524
rect 22235 34493 22247 34496
rect 22189 34487 22247 34493
rect 23492 34456 23520 34496
rect 23934 34484 23940 34536
rect 23992 34524 23998 34536
rect 24949 34527 25007 34533
rect 24949 34524 24961 34527
rect 23992 34496 24961 34524
rect 23992 34484 23998 34496
rect 24949 34493 24961 34496
rect 24995 34524 25007 34527
rect 26050 34524 26056 34536
rect 24995 34496 26056 34524
rect 24995 34493 25007 34496
rect 24949 34487 25007 34493
rect 26050 34484 26056 34496
rect 26108 34484 26114 34536
rect 29181 34527 29239 34533
rect 29181 34493 29193 34527
rect 29227 34524 29239 34527
rect 29454 34524 29460 34536
rect 29227 34496 29460 34524
rect 29227 34493 29239 34496
rect 29181 34487 29239 34493
rect 29454 34484 29460 34496
rect 29512 34484 29518 34536
rect 30009 34527 30067 34533
rect 30009 34493 30021 34527
rect 30055 34524 30067 34527
rect 30374 34524 30380 34536
rect 30055 34496 30380 34524
rect 30055 34493 30067 34496
rect 30009 34487 30067 34493
rect 30374 34484 30380 34496
rect 30432 34484 30438 34536
rect 30466 34484 30472 34536
rect 30524 34524 30530 34536
rect 30852 34524 30880 34555
rect 31202 34552 31208 34564
rect 31260 34552 31266 34604
rect 31478 34592 31484 34604
rect 31439 34564 31484 34592
rect 31478 34552 31484 34564
rect 31536 34552 31542 34604
rect 31662 34592 31668 34604
rect 31623 34564 31668 34592
rect 31662 34552 31668 34564
rect 31720 34552 31726 34604
rect 30524 34496 30880 34524
rect 30524 34484 30530 34496
rect 24854 34456 24860 34468
rect 22020 34428 22094 34456
rect 23492 34428 24860 34456
rect 16080 34416 16086 34428
rect 10505 34391 10563 34397
rect 10505 34357 10517 34391
rect 10551 34388 10563 34391
rect 10686 34388 10692 34400
rect 10551 34360 10692 34388
rect 10551 34357 10563 34360
rect 10505 34351 10563 34357
rect 10686 34348 10692 34360
rect 10744 34348 10750 34400
rect 14479 34391 14537 34397
rect 14479 34357 14491 34391
rect 14525 34388 14537 34391
rect 16114 34388 16120 34400
rect 14525 34360 16120 34388
rect 14525 34357 14537 34360
rect 14479 34351 14537 34357
rect 16114 34348 16120 34360
rect 16172 34348 16178 34400
rect 17497 34391 17555 34397
rect 17497 34357 17509 34391
rect 17543 34388 17555 34391
rect 17862 34388 17868 34400
rect 17543 34360 17868 34388
rect 17543 34357 17555 34360
rect 17497 34351 17555 34357
rect 17862 34348 17868 34360
rect 17920 34348 17926 34400
rect 18230 34348 18236 34400
rect 18288 34388 18294 34400
rect 19686 34391 19744 34397
rect 19686 34388 19698 34391
rect 18288 34360 19698 34388
rect 18288 34348 18294 34360
rect 19686 34357 19698 34360
rect 19732 34357 19744 34391
rect 22066 34388 22094 34428
rect 24854 34416 24860 34428
rect 24912 34416 24918 34468
rect 30282 34456 30288 34468
rect 30243 34428 30288 34456
rect 30282 34416 30288 34428
rect 30340 34416 30346 34468
rect 33594 34456 33600 34468
rect 33555 34428 33600 34456
rect 33594 34416 33600 34428
rect 33652 34416 33658 34468
rect 22186 34388 22192 34400
rect 22066 34360 22192 34388
rect 19686 34351 19744 34357
rect 22186 34348 22192 34360
rect 22244 34348 22250 34400
rect 24394 34388 24400 34400
rect 24355 34360 24400 34388
rect 24394 34348 24400 34360
rect 24452 34348 24458 34400
rect 26234 34388 26240 34400
rect 26195 34360 26240 34388
rect 26234 34348 26240 34360
rect 26292 34348 26298 34400
rect 27890 34348 27896 34400
rect 27948 34388 27954 34400
rect 27985 34391 28043 34397
rect 27985 34388 27997 34391
rect 27948 34360 27997 34388
rect 27948 34348 27954 34360
rect 27985 34357 27997 34360
rect 28031 34388 28043 34391
rect 28626 34388 28632 34400
rect 28031 34360 28632 34388
rect 28031 34357 28043 34360
rect 27985 34351 28043 34357
rect 28626 34348 28632 34360
rect 28684 34348 28690 34400
rect 1104 34298 37628 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 37628 34298
rect 1104 34224 37628 34246
rect 12158 34144 12164 34196
rect 12216 34184 12222 34196
rect 12621 34187 12679 34193
rect 12621 34184 12633 34187
rect 12216 34156 12633 34184
rect 12216 34144 12222 34156
rect 12621 34153 12633 34156
rect 12667 34153 12679 34187
rect 12621 34147 12679 34153
rect 15013 34187 15071 34193
rect 15013 34153 15025 34187
rect 15059 34184 15071 34187
rect 15286 34184 15292 34196
rect 15059 34156 15292 34184
rect 15059 34153 15071 34156
rect 15013 34147 15071 34153
rect 15286 34144 15292 34156
rect 15344 34144 15350 34196
rect 18230 34184 18236 34196
rect 18191 34156 18236 34184
rect 18230 34144 18236 34156
rect 18288 34144 18294 34196
rect 20806 34184 20812 34196
rect 18340 34156 19656 34184
rect 20767 34156 20812 34184
rect 17034 34076 17040 34128
rect 17092 34116 17098 34128
rect 18340 34116 18368 34156
rect 17092 34088 18368 34116
rect 19521 34119 19579 34125
rect 17092 34076 17098 34088
rect 19521 34085 19533 34119
rect 19567 34085 19579 34119
rect 19628 34116 19656 34156
rect 20806 34144 20812 34156
rect 20864 34144 20870 34196
rect 26694 34184 26700 34196
rect 26655 34156 26700 34184
rect 26694 34144 26700 34156
rect 26752 34144 26758 34196
rect 27706 34144 27712 34196
rect 27764 34184 27770 34196
rect 27801 34187 27859 34193
rect 27801 34184 27813 34187
rect 27764 34156 27813 34184
rect 27764 34144 27770 34156
rect 27801 34153 27813 34156
rect 27847 34153 27859 34187
rect 33134 34184 33140 34196
rect 33095 34156 33140 34184
rect 27801 34147 27859 34153
rect 33134 34144 33140 34156
rect 33192 34144 33198 34196
rect 28258 34116 28264 34128
rect 19628 34088 20944 34116
rect 19521 34079 19579 34085
rect 8018 34008 8024 34060
rect 8076 34048 8082 34060
rect 8389 34051 8447 34057
rect 8389 34048 8401 34051
rect 8076 34020 8401 34048
rect 8076 34008 8082 34020
rect 8389 34017 8401 34020
rect 8435 34017 8447 34051
rect 8389 34011 8447 34017
rect 9490 34008 9496 34060
rect 9548 34048 9554 34060
rect 9585 34051 9643 34057
rect 9585 34048 9597 34051
rect 9548 34020 9597 34048
rect 9548 34008 9554 34020
rect 9585 34017 9597 34020
rect 9631 34017 9643 34051
rect 9585 34011 9643 34017
rect 9674 34008 9680 34060
rect 9732 34048 9738 34060
rect 10686 34048 10692 34060
rect 9732 34020 9777 34048
rect 10647 34020 10692 34048
rect 9732 34008 9738 34020
rect 10686 34008 10692 34020
rect 10744 34008 10750 34060
rect 12526 34008 12532 34060
rect 12584 34048 12590 34060
rect 13173 34051 13231 34057
rect 13173 34048 13185 34051
rect 12584 34020 13185 34048
rect 12584 34008 12590 34020
rect 13173 34017 13185 34020
rect 13219 34017 13231 34051
rect 13173 34011 13231 34017
rect 14182 34008 14188 34060
rect 14240 34048 14246 34060
rect 14369 34051 14427 34057
rect 14369 34048 14381 34051
rect 14240 34020 14381 34048
rect 14240 34008 14246 34020
rect 14369 34017 14381 34020
rect 14415 34048 14427 34051
rect 14642 34048 14648 34060
rect 14415 34020 14648 34048
rect 14415 34017 14427 34020
rect 14369 34011 14427 34017
rect 14642 34008 14648 34020
rect 14700 34008 14706 34060
rect 16022 34008 16028 34060
rect 16080 34048 16086 34060
rect 16117 34051 16175 34057
rect 16117 34048 16129 34051
rect 16080 34020 16129 34048
rect 16080 34008 16086 34020
rect 16117 34017 16129 34020
rect 16163 34017 16175 34051
rect 16117 34011 16175 34017
rect 8202 33940 8208 33992
rect 8260 33980 8266 33992
rect 9766 33980 9772 33992
rect 8260 33952 9772 33980
rect 8260 33940 8266 33952
rect 9766 33940 9772 33952
rect 9824 33980 9830 33992
rect 10410 33980 10416 33992
rect 9824 33952 10416 33980
rect 9824 33940 9830 33952
rect 10410 33940 10416 33952
rect 10468 33940 10474 33992
rect 13081 33983 13139 33989
rect 13081 33980 13093 33983
rect 12176 33952 13093 33980
rect 8478 33912 8484 33924
rect 8220 33884 8484 33912
rect 7374 33804 7380 33856
rect 7432 33844 7438 33856
rect 8220 33853 8248 33884
rect 8478 33872 8484 33884
rect 8536 33872 8542 33924
rect 9582 33912 9588 33924
rect 8956 33884 9588 33912
rect 7837 33847 7895 33853
rect 7837 33844 7849 33847
rect 7432 33816 7849 33844
rect 7432 33804 7438 33816
rect 7837 33813 7849 33816
rect 7883 33813 7895 33847
rect 7837 33807 7895 33813
rect 8205 33847 8263 33853
rect 8205 33813 8217 33847
rect 8251 33813 8263 33847
rect 8205 33807 8263 33813
rect 8297 33847 8355 33853
rect 8297 33813 8309 33847
rect 8343 33844 8355 33847
rect 8956 33844 8984 33884
rect 9582 33872 9588 33884
rect 9640 33872 9646 33924
rect 11146 33872 11152 33924
rect 11204 33872 11210 33924
rect 12176 33856 12204 33952
rect 13081 33949 13093 33952
rect 13127 33949 13139 33983
rect 15930 33980 15936 33992
rect 15891 33952 15936 33980
rect 13081 33943 13139 33949
rect 15930 33940 15936 33952
rect 15988 33940 15994 33992
rect 16761 33983 16819 33989
rect 16761 33949 16773 33983
rect 16807 33980 16819 33983
rect 17052 33980 17080 34076
rect 19334 34048 19340 34060
rect 18064 34020 19340 34048
rect 17402 33980 17408 33992
rect 16807 33952 17080 33980
rect 17363 33952 17408 33980
rect 16807 33949 16819 33952
rect 16761 33943 16819 33949
rect 17402 33940 17408 33952
rect 17460 33940 17466 33992
rect 18064 33989 18092 34020
rect 19334 34008 19340 34020
rect 19392 34008 19398 34060
rect 18049 33983 18107 33989
rect 18049 33949 18061 33983
rect 18095 33949 18107 33983
rect 18049 33943 18107 33949
rect 18693 33983 18751 33989
rect 18693 33949 18705 33983
rect 18739 33980 18751 33983
rect 19536 33980 19564 34079
rect 19978 34008 19984 34060
rect 20036 34048 20042 34060
rect 20073 34051 20131 34057
rect 20073 34048 20085 34051
rect 20036 34020 20085 34048
rect 20036 34008 20042 34020
rect 20073 34017 20085 34020
rect 20119 34017 20131 34051
rect 20073 34011 20131 34017
rect 20916 33992 20944 34088
rect 28000 34088 28264 34116
rect 23382 34048 23388 34060
rect 23343 34020 23388 34048
rect 23382 34008 23388 34020
rect 23440 34008 23446 34060
rect 24854 34008 24860 34060
rect 24912 34048 24918 34060
rect 24949 34051 25007 34057
rect 24949 34048 24961 34051
rect 24912 34020 24961 34048
rect 24912 34008 24918 34020
rect 24949 34017 24961 34020
rect 24995 34017 25007 34051
rect 24949 34011 25007 34017
rect 25225 34051 25283 34057
rect 25225 34017 25237 34051
rect 25271 34048 25283 34051
rect 26234 34048 26240 34060
rect 25271 34020 26240 34048
rect 25271 34017 25283 34020
rect 25225 34011 25283 34017
rect 26234 34008 26240 34020
rect 26292 34008 26298 34060
rect 20898 33980 20904 33992
rect 18739 33952 19564 33980
rect 20859 33952 20904 33980
rect 18739 33949 18751 33952
rect 18693 33943 18751 33949
rect 20898 33940 20904 33952
rect 20956 33980 20962 33992
rect 21266 33980 21272 33992
rect 20956 33952 21272 33980
rect 20956 33940 20962 33952
rect 21266 33940 21272 33952
rect 21324 33940 21330 33992
rect 21358 33940 21364 33992
rect 21416 33980 21422 33992
rect 22189 33983 22247 33989
rect 22189 33980 22201 33983
rect 21416 33952 22201 33980
rect 21416 33940 21422 33952
rect 22189 33949 22201 33952
rect 22235 33949 22247 33983
rect 22189 33943 22247 33949
rect 23201 33983 23259 33989
rect 23201 33949 23213 33983
rect 23247 33980 23259 33983
rect 24394 33980 24400 33992
rect 23247 33952 24400 33980
rect 23247 33949 23259 33952
rect 23201 33943 23259 33949
rect 24394 33940 24400 33952
rect 24452 33940 24458 33992
rect 28000 33989 28028 34088
rect 28258 34076 28264 34088
rect 28316 34076 28322 34128
rect 27985 33983 28043 33989
rect 27985 33949 27997 33983
rect 28031 33949 28043 33983
rect 27985 33943 28043 33949
rect 28077 33983 28135 33989
rect 28077 33949 28089 33983
rect 28123 33949 28135 33983
rect 28077 33943 28135 33949
rect 14553 33915 14611 33921
rect 14553 33912 14565 33915
rect 13004 33884 14565 33912
rect 9122 33844 9128 33856
rect 8343 33816 8984 33844
rect 9083 33816 9128 33844
rect 8343 33813 8355 33816
rect 8297 33807 8355 33813
rect 9122 33804 9128 33816
rect 9180 33804 9186 33856
rect 9490 33844 9496 33856
rect 9451 33816 9496 33844
rect 9490 33804 9496 33816
rect 9548 33804 9554 33856
rect 11974 33804 11980 33856
rect 12032 33844 12038 33856
rect 12158 33844 12164 33856
rect 12032 33816 12164 33844
rect 12032 33804 12038 33816
rect 12158 33804 12164 33816
rect 12216 33804 12222 33856
rect 12894 33804 12900 33856
rect 12952 33844 12958 33856
rect 13004 33853 13032 33884
rect 14553 33881 14565 33884
rect 14599 33881 14611 33915
rect 14553 33875 14611 33881
rect 19058 33872 19064 33924
rect 19116 33912 19122 33924
rect 19981 33915 20039 33921
rect 19981 33912 19993 33915
rect 19116 33884 19993 33912
rect 19116 33872 19122 33884
rect 19981 33881 19993 33884
rect 20027 33881 20039 33915
rect 26602 33912 26608 33924
rect 26450 33884 26608 33912
rect 19981 33875 20039 33881
rect 26602 33872 26608 33884
rect 26660 33872 26666 33924
rect 28092 33912 28120 33943
rect 28166 33940 28172 33992
rect 28224 33980 28230 33992
rect 28261 33983 28319 33989
rect 28261 33980 28273 33983
rect 28224 33952 28273 33980
rect 28224 33940 28230 33952
rect 28261 33949 28273 33952
rect 28307 33949 28319 33983
rect 28261 33943 28319 33949
rect 28353 33983 28411 33989
rect 28353 33949 28365 33983
rect 28399 33980 28411 33983
rect 28534 33980 28540 33992
rect 28399 33952 28540 33980
rect 28399 33949 28411 33952
rect 28353 33943 28411 33949
rect 28534 33940 28540 33952
rect 28592 33940 28598 33992
rect 28626 33940 28632 33992
rect 28684 33980 28690 33992
rect 29917 33983 29975 33989
rect 29917 33980 29929 33983
rect 28684 33952 29929 33980
rect 28684 33940 28690 33952
rect 29917 33949 29929 33952
rect 29963 33980 29975 33983
rect 30466 33980 30472 33992
rect 29963 33952 30472 33980
rect 29963 33949 29975 33952
rect 29917 33943 29975 33949
rect 30466 33940 30472 33952
rect 30524 33940 30530 33992
rect 32585 33983 32643 33989
rect 32585 33949 32597 33983
rect 32631 33980 32643 33983
rect 32766 33980 32772 33992
rect 32631 33952 32772 33980
rect 32631 33949 32643 33952
rect 32585 33943 32643 33949
rect 32766 33940 32772 33952
rect 32824 33940 32830 33992
rect 33229 33983 33287 33989
rect 33229 33949 33241 33983
rect 33275 33980 33287 33983
rect 33502 33980 33508 33992
rect 33275 33952 33508 33980
rect 33275 33949 33287 33952
rect 33229 33943 33287 33949
rect 33502 33940 33508 33952
rect 33560 33940 33566 33992
rect 28442 33912 28448 33924
rect 28092 33884 28448 33912
rect 28442 33872 28448 33884
rect 28500 33872 28506 33924
rect 32309 33915 32367 33921
rect 31878 33884 32260 33912
rect 12989 33847 13047 33853
rect 12989 33844 13001 33847
rect 12952 33816 13001 33844
rect 12952 33804 12958 33816
rect 12989 33813 13001 33816
rect 13035 33813 13047 33847
rect 12989 33807 13047 33813
rect 13906 33804 13912 33856
rect 13964 33844 13970 33856
rect 14645 33847 14703 33853
rect 14645 33844 14657 33847
rect 13964 33816 14657 33844
rect 13964 33804 13970 33816
rect 14645 33813 14657 33816
rect 14691 33813 14703 33847
rect 15562 33844 15568 33856
rect 15523 33816 15568 33844
rect 14645 33807 14703 33813
rect 15562 33804 15568 33816
rect 15620 33804 15626 33856
rect 16025 33847 16083 33853
rect 16025 33813 16037 33847
rect 16071 33844 16083 33847
rect 16574 33844 16580 33856
rect 16071 33816 16580 33844
rect 16071 33813 16083 33816
rect 16025 33807 16083 33813
rect 16574 33804 16580 33816
rect 16632 33804 16638 33856
rect 16850 33844 16856 33856
rect 16811 33816 16856 33844
rect 16850 33804 16856 33816
rect 16908 33804 16914 33856
rect 17586 33844 17592 33856
rect 17547 33816 17592 33844
rect 17586 33804 17592 33816
rect 17644 33804 17650 33856
rect 18874 33844 18880 33856
rect 18835 33816 18880 33844
rect 18874 33804 18880 33816
rect 18932 33804 18938 33856
rect 19794 33804 19800 33856
rect 19852 33844 19858 33856
rect 19889 33847 19947 33853
rect 19889 33844 19901 33847
rect 19852 33816 19901 33844
rect 19852 33804 19858 33816
rect 19889 33813 19901 33816
rect 19935 33813 19947 33847
rect 22278 33844 22284 33856
rect 22239 33816 22284 33844
rect 19889 33807 19947 33813
rect 22278 33804 22284 33816
rect 22336 33804 22342 33856
rect 22830 33844 22836 33856
rect 22791 33816 22836 33844
rect 22830 33804 22836 33816
rect 22888 33804 22894 33856
rect 23293 33847 23351 33853
rect 23293 33813 23305 33847
rect 23339 33844 23351 33847
rect 23842 33844 23848 33856
rect 23339 33816 23848 33844
rect 23339 33813 23351 33816
rect 23293 33807 23351 33813
rect 23842 33804 23848 33816
rect 23900 33804 23906 33856
rect 28534 33804 28540 33856
rect 28592 33844 28598 33856
rect 29825 33847 29883 33853
rect 29825 33844 29837 33847
rect 28592 33816 29837 33844
rect 28592 33804 28598 33816
rect 29825 33813 29837 33816
rect 29871 33844 29883 33847
rect 29914 33844 29920 33856
rect 29871 33816 29920 33844
rect 29871 33813 29883 33816
rect 29825 33807 29883 33813
rect 29914 33804 29920 33816
rect 29972 33804 29978 33856
rect 30098 33804 30104 33856
rect 30156 33844 30162 33856
rect 30837 33847 30895 33853
rect 30837 33844 30849 33847
rect 30156 33816 30849 33844
rect 30156 33804 30162 33816
rect 30837 33813 30849 33816
rect 30883 33813 30895 33847
rect 32232 33844 32260 33884
rect 32309 33881 32321 33915
rect 32355 33912 32367 33915
rect 32398 33912 32404 33924
rect 32355 33884 32404 33912
rect 32355 33881 32367 33884
rect 32309 33875 32367 33881
rect 32398 33872 32404 33884
rect 32456 33872 32462 33924
rect 33042 33844 33048 33856
rect 32232 33816 33048 33844
rect 30837 33807 30895 33813
rect 33042 33804 33048 33816
rect 33100 33804 33106 33856
rect 1104 33754 37628 33776
rect 1104 33702 4874 33754
rect 4926 33702 4938 33754
rect 4990 33702 5002 33754
rect 5054 33702 5066 33754
rect 5118 33702 5130 33754
rect 5182 33702 35594 33754
rect 35646 33702 35658 33754
rect 35710 33702 35722 33754
rect 35774 33702 35786 33754
rect 35838 33702 35850 33754
rect 35902 33702 37628 33754
rect 1104 33680 37628 33702
rect 9582 33640 9588 33652
rect 9543 33612 9588 33640
rect 9582 33600 9588 33612
rect 9640 33600 9646 33652
rect 10502 33600 10508 33652
rect 10560 33640 10566 33652
rect 10781 33643 10839 33649
rect 10781 33640 10793 33643
rect 10560 33612 10793 33640
rect 10560 33600 10566 33612
rect 10781 33609 10793 33612
rect 10827 33609 10839 33643
rect 10781 33603 10839 33609
rect 15565 33643 15623 33649
rect 15565 33609 15577 33643
rect 15611 33609 15623 33643
rect 15565 33603 15623 33609
rect 15933 33643 15991 33649
rect 15933 33609 15945 33643
rect 15979 33640 15991 33643
rect 16574 33640 16580 33652
rect 15979 33612 16580 33640
rect 15979 33609 15991 33612
rect 15933 33603 15991 33609
rect 6914 33532 6920 33584
rect 6972 33572 6978 33584
rect 8202 33572 8208 33584
rect 6972 33544 8208 33572
rect 6972 33532 6978 33544
rect 7374 33504 7380 33516
rect 7335 33476 7380 33504
rect 7374 33464 7380 33476
rect 7432 33464 7438 33516
rect 7852 33513 7880 33544
rect 8202 33532 8208 33544
rect 8260 33532 8266 33584
rect 8386 33532 8392 33584
rect 8444 33572 8450 33584
rect 8444 33544 8602 33572
rect 8444 33532 8450 33544
rect 10134 33532 10140 33584
rect 10192 33572 10198 33584
rect 10413 33575 10471 33581
rect 10413 33572 10425 33575
rect 10192 33544 10425 33572
rect 10192 33532 10198 33544
rect 10413 33541 10425 33544
rect 10459 33541 10471 33575
rect 10413 33535 10471 33541
rect 11790 33532 11796 33584
rect 11848 33572 11854 33584
rect 12529 33575 12587 33581
rect 12529 33572 12541 33575
rect 11848 33544 12541 33572
rect 11848 33532 11854 33544
rect 12529 33541 12541 33544
rect 12575 33541 12587 33575
rect 12529 33535 12587 33541
rect 12986 33532 12992 33584
rect 13044 33532 13050 33584
rect 7837 33507 7895 33513
rect 7837 33473 7849 33507
rect 7883 33473 7895 33507
rect 7837 33467 7895 33473
rect 10042 33464 10048 33516
rect 10100 33504 10106 33516
rect 10321 33507 10379 33513
rect 10321 33504 10333 33507
rect 10100 33476 10333 33504
rect 10100 33464 10106 33476
rect 10321 33473 10333 33476
rect 10367 33473 10379 33507
rect 10321 33467 10379 33473
rect 14921 33507 14979 33513
rect 14921 33473 14933 33507
rect 14967 33504 14979 33507
rect 15580 33504 15608 33603
rect 16574 33600 16580 33612
rect 16632 33640 16638 33652
rect 17494 33640 17500 33652
rect 16632 33612 17500 33640
rect 16632 33600 16638 33612
rect 17494 33600 17500 33612
rect 17552 33600 17558 33652
rect 18414 33600 18420 33652
rect 18472 33640 18478 33652
rect 19058 33640 19064 33652
rect 18472 33612 19064 33640
rect 18472 33600 18478 33612
rect 19058 33600 19064 33612
rect 19116 33600 19122 33652
rect 22094 33640 22100 33652
rect 22066 33600 22100 33640
rect 22152 33600 22158 33652
rect 30098 33600 30104 33652
rect 30156 33640 30162 33652
rect 32398 33640 32404 33652
rect 30156 33612 30880 33640
rect 32359 33612 32404 33640
rect 30156 33600 30162 33612
rect 17586 33572 17592 33584
rect 17547 33544 17592 33572
rect 17586 33532 17592 33544
rect 17644 33532 17650 33584
rect 17862 33532 17868 33584
rect 17920 33572 17926 33584
rect 17920 33544 18078 33572
rect 17920 33532 17926 33544
rect 19426 33532 19432 33584
rect 19484 33572 19490 33584
rect 19613 33575 19671 33581
rect 19613 33572 19625 33575
rect 19484 33544 19625 33572
rect 19484 33532 19490 33544
rect 19613 33541 19625 33544
rect 19659 33541 19671 33575
rect 22066 33572 22094 33600
rect 19613 33535 19671 33541
rect 22020 33544 22094 33572
rect 17126 33504 17132 33516
rect 14967 33476 15608 33504
rect 16224 33476 17132 33504
rect 14967 33473 14979 33476
rect 14921 33467 14979 33473
rect 16224 33448 16252 33476
rect 17126 33464 17132 33476
rect 17184 33464 17190 33516
rect 20441 33507 20499 33513
rect 20441 33473 20453 33507
rect 20487 33504 20499 33507
rect 20714 33504 20720 33516
rect 20487 33476 20720 33504
rect 20487 33473 20499 33476
rect 20441 33467 20499 33473
rect 20714 33464 20720 33476
rect 20772 33504 20778 33516
rect 21818 33504 21824 33516
rect 20772 33476 21824 33504
rect 20772 33464 20778 33476
rect 21818 33464 21824 33476
rect 21876 33464 21882 33516
rect 22020 33513 22048 33544
rect 22278 33532 22284 33584
rect 22336 33572 22342 33584
rect 30653 33575 30711 33581
rect 30653 33572 30665 33575
rect 22336 33544 22770 33572
rect 29380 33544 30665 33572
rect 22336 33532 22342 33544
rect 22005 33507 22063 33513
rect 22005 33473 22017 33507
rect 22051 33473 22063 33507
rect 24210 33504 24216 33516
rect 24171 33476 24216 33504
rect 22005 33467 22063 33473
rect 24210 33464 24216 33476
rect 24268 33464 24274 33516
rect 24854 33504 24860 33516
rect 24815 33476 24860 33504
rect 24854 33464 24860 33476
rect 24912 33464 24918 33516
rect 26234 33464 26240 33516
rect 26292 33464 26298 33516
rect 29380 33513 29408 33544
rect 30653 33541 30665 33544
rect 30699 33541 30711 33575
rect 30653 33535 30711 33541
rect 29365 33507 29423 33513
rect 29365 33473 29377 33507
rect 29411 33473 29423 33507
rect 29365 33467 29423 33473
rect 30006 33464 30012 33516
rect 30064 33504 30070 33516
rect 30561 33507 30619 33513
rect 30561 33504 30573 33507
rect 30064 33476 30573 33504
rect 30064 33464 30070 33476
rect 30561 33473 30573 33476
rect 30607 33473 30619 33507
rect 30561 33467 30619 33473
rect 30745 33507 30803 33513
rect 30745 33473 30757 33507
rect 30791 33473 30803 33507
rect 30852 33504 30880 33612
rect 32398 33600 32404 33612
rect 32456 33600 32462 33652
rect 33042 33640 33048 33652
rect 33003 33612 33048 33640
rect 33042 33600 33048 33612
rect 33100 33600 33106 33652
rect 31205 33507 31263 33513
rect 31205 33504 31217 33507
rect 30852 33476 31217 33504
rect 30745 33467 30803 33473
rect 31205 33473 31217 33476
rect 31251 33473 31263 33507
rect 31386 33504 31392 33516
rect 31347 33476 31392 33504
rect 31205 33467 31263 33473
rect 8110 33436 8116 33448
rect 8071 33408 8116 33436
rect 8110 33396 8116 33408
rect 8168 33396 8174 33448
rect 10229 33439 10287 33445
rect 10229 33405 10241 33439
rect 10275 33436 10287 33439
rect 10962 33436 10968 33448
rect 10275 33408 10968 33436
rect 10275 33405 10287 33408
rect 10229 33399 10287 33405
rect 10962 33396 10968 33408
rect 11020 33436 11026 33448
rect 12250 33436 12256 33448
rect 11020 33408 12112 33436
rect 12211 33408 12256 33436
rect 11020 33396 11026 33408
rect 7006 33260 7012 33312
rect 7064 33300 7070 33312
rect 7193 33303 7251 33309
rect 7193 33300 7205 33303
rect 7064 33272 7205 33300
rect 7064 33260 7070 33272
rect 7193 33269 7205 33272
rect 7239 33269 7251 33303
rect 12084 33300 12112 33408
rect 12250 33396 12256 33408
rect 12308 33396 12314 33448
rect 12894 33396 12900 33448
rect 12952 33436 12958 33448
rect 14001 33439 14059 33445
rect 14001 33436 14013 33439
rect 12952 33408 14013 33436
rect 12952 33396 12958 33408
rect 14001 33405 14013 33408
rect 14047 33405 14059 33439
rect 16022 33436 16028 33448
rect 15983 33408 16028 33436
rect 14001 33399 14059 33405
rect 16022 33396 16028 33408
rect 16080 33396 16086 33448
rect 16206 33436 16212 33448
rect 16167 33408 16212 33436
rect 16206 33396 16212 33408
rect 16264 33396 16270 33448
rect 16666 33396 16672 33448
rect 16724 33436 16730 33448
rect 17313 33439 17371 33445
rect 17313 33436 17325 33439
rect 16724 33408 17325 33436
rect 16724 33396 16730 33408
rect 17313 33405 17325 33408
rect 17359 33405 17371 33439
rect 22278 33436 22284 33448
rect 22239 33408 22284 33436
rect 17313 33399 17371 33405
rect 22278 33396 22284 33408
rect 22336 33396 22342 33448
rect 25133 33439 25191 33445
rect 25133 33436 25145 33439
rect 24412 33408 25145 33436
rect 24412 33377 24440 33408
rect 25133 33405 25145 33408
rect 25179 33405 25191 33439
rect 25133 33399 25191 33405
rect 27706 33396 27712 33448
rect 27764 33436 27770 33448
rect 28077 33439 28135 33445
rect 28077 33436 28089 33439
rect 27764 33408 28089 33436
rect 27764 33396 27770 33408
rect 28077 33405 28089 33408
rect 28123 33405 28135 33439
rect 28077 33399 28135 33405
rect 28537 33439 28595 33445
rect 28537 33405 28549 33439
rect 28583 33436 28595 33439
rect 28583 33408 29132 33436
rect 28583 33405 28595 33408
rect 28537 33399 28595 33405
rect 24397 33371 24455 33377
rect 24397 33337 24409 33371
rect 24443 33337 24455 33371
rect 24397 33331 24455 33337
rect 26694 33328 26700 33380
rect 26752 33368 26758 33380
rect 28353 33371 28411 33377
rect 28353 33368 28365 33371
rect 26752 33340 28365 33368
rect 26752 33328 26758 33340
rect 28353 33337 28365 33340
rect 28399 33337 28411 33371
rect 28994 33368 29000 33380
rect 28955 33340 29000 33368
rect 28353 33331 28411 33337
rect 28994 33328 29000 33340
rect 29052 33328 29058 33380
rect 29104 33368 29132 33408
rect 29178 33396 29184 33448
rect 29236 33436 29242 33448
rect 29236 33408 29281 33436
rect 29236 33396 29242 33408
rect 29914 33396 29920 33448
rect 29972 33436 29978 33448
rect 30760 33436 30788 33467
rect 31386 33464 31392 33476
rect 31444 33464 31450 33516
rect 32309 33507 32367 33513
rect 32309 33504 32321 33507
rect 31726 33476 32321 33504
rect 29972 33408 30788 33436
rect 31297 33439 31355 33445
rect 29972 33396 29978 33408
rect 31297 33405 31309 33439
rect 31343 33436 31355 33439
rect 31726 33436 31754 33476
rect 32309 33473 32321 33476
rect 32355 33473 32367 33507
rect 32309 33467 32367 33473
rect 32493 33507 32551 33513
rect 32493 33473 32505 33507
rect 32539 33473 32551 33507
rect 32493 33467 32551 33473
rect 33137 33507 33195 33513
rect 33137 33473 33149 33507
rect 33183 33504 33195 33507
rect 33502 33504 33508 33516
rect 33183 33476 33508 33504
rect 33183 33473 33195 33476
rect 33137 33467 33195 33473
rect 31343 33408 31754 33436
rect 31343 33405 31355 33408
rect 31297 33399 31355 33405
rect 29273 33371 29331 33377
rect 29273 33368 29285 33371
rect 29104 33340 29285 33368
rect 29273 33337 29285 33340
rect 29319 33368 29331 33371
rect 29638 33368 29644 33380
rect 29319 33340 29644 33368
rect 29319 33337 29331 33340
rect 29273 33331 29331 33337
rect 29638 33328 29644 33340
rect 29696 33328 29702 33380
rect 30374 33328 30380 33380
rect 30432 33368 30438 33380
rect 32508 33368 32536 33467
rect 33502 33464 33508 33476
rect 33560 33504 33566 33516
rect 33778 33504 33784 33516
rect 33560 33476 33784 33504
rect 33560 33464 33566 33476
rect 33778 33464 33784 33476
rect 33836 33464 33842 33516
rect 30432 33340 32536 33368
rect 30432 33328 30438 33340
rect 14182 33300 14188 33312
rect 12084 33272 14188 33300
rect 7193 33263 7251 33269
rect 14182 33260 14188 33272
rect 14240 33260 14246 33312
rect 15102 33300 15108 33312
rect 15063 33272 15108 33300
rect 15102 33260 15108 33272
rect 15160 33260 15166 33312
rect 23753 33303 23811 33309
rect 23753 33269 23765 33303
rect 23799 33300 23811 33303
rect 23842 33300 23848 33312
rect 23799 33272 23848 33300
rect 23799 33269 23811 33272
rect 23753 33263 23811 33269
rect 23842 33260 23848 33272
rect 23900 33260 23906 33312
rect 24946 33260 24952 33312
rect 25004 33300 25010 33312
rect 26605 33303 26663 33309
rect 26605 33300 26617 33303
rect 25004 33272 26617 33300
rect 25004 33260 25010 33272
rect 26605 33269 26617 33272
rect 26651 33300 26663 33303
rect 27522 33300 27528 33312
rect 26651 33272 27528 33300
rect 26651 33269 26663 33272
rect 26605 33263 26663 33269
rect 27522 33260 27528 33272
rect 27580 33260 27586 33312
rect 29178 33300 29184 33312
rect 29139 33272 29184 33300
rect 29178 33260 29184 33272
rect 29236 33260 29242 33312
rect 1104 33210 37628 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 37628 33210
rect 1104 33136 37628 33158
rect 8478 33096 8484 33108
rect 8439 33068 8484 33096
rect 8478 33056 8484 33068
rect 8536 33056 8542 33108
rect 9490 33056 9496 33108
rect 9548 33096 9554 33108
rect 9585 33099 9643 33105
rect 9585 33096 9597 33099
rect 9548 33068 9597 33096
rect 9548 33056 9554 33068
rect 9585 33065 9597 33068
rect 9631 33065 9643 33099
rect 9585 33059 9643 33065
rect 12066 33056 12072 33108
rect 12124 33096 12130 33108
rect 12345 33099 12403 33105
rect 12345 33096 12357 33099
rect 12124 33068 12357 33096
rect 12124 33056 12130 33068
rect 12345 33065 12357 33068
rect 12391 33065 12403 33099
rect 12345 33059 12403 33065
rect 14274 33056 14280 33108
rect 14332 33096 14338 33108
rect 14645 33099 14703 33105
rect 14645 33096 14657 33099
rect 14332 33068 14657 33096
rect 14332 33056 14338 33068
rect 14645 33065 14657 33068
rect 14691 33065 14703 33099
rect 14645 33059 14703 33065
rect 15102 33056 15108 33108
rect 15160 33096 15166 33108
rect 16098 33099 16156 33105
rect 16098 33096 16110 33099
rect 15160 33068 16110 33096
rect 15160 33056 15166 33068
rect 16098 33065 16110 33068
rect 16144 33065 16156 33099
rect 16098 33059 16156 33065
rect 17402 33056 17408 33108
rect 17460 33096 17466 33108
rect 18141 33099 18199 33105
rect 18141 33096 18153 33099
rect 17460 33068 18153 33096
rect 17460 33056 17466 33068
rect 18141 33065 18153 33068
rect 18187 33065 18199 33099
rect 19518 33096 19524 33108
rect 18141 33059 18199 33065
rect 18708 33068 19524 33096
rect 7006 32960 7012 32972
rect 6967 32932 7012 32960
rect 7006 32920 7012 32932
rect 7064 32920 7070 32972
rect 8496 32960 8524 33056
rect 12618 33028 12624 33040
rect 11716 33000 12624 33028
rect 10042 32960 10048 32972
rect 8496 32932 10048 32960
rect 10042 32920 10048 32932
rect 10100 32920 10106 32972
rect 10229 32963 10287 32969
rect 10229 32929 10241 32963
rect 10275 32960 10287 32963
rect 10318 32960 10324 32972
rect 10275 32932 10324 32960
rect 10275 32929 10287 32932
rect 10229 32923 10287 32929
rect 6454 32852 6460 32904
rect 6512 32892 6518 32904
rect 6730 32892 6736 32904
rect 6512 32864 6736 32892
rect 6512 32852 6518 32864
rect 6730 32852 6736 32864
rect 6788 32852 6794 32904
rect 9674 32852 9680 32904
rect 9732 32892 9738 32904
rect 10244 32892 10272 32923
rect 10318 32920 10324 32932
rect 10376 32960 10382 32972
rect 11716 32969 11744 33000
rect 12618 32988 12624 33000
rect 12676 32988 12682 33040
rect 15562 33028 15568 33040
rect 15120 33000 15568 33028
rect 11701 32963 11759 32969
rect 11701 32960 11713 32963
rect 10376 32932 11713 32960
rect 10376 32920 10382 32932
rect 11701 32929 11713 32932
rect 11747 32929 11759 32963
rect 11701 32923 11759 32929
rect 11885 32963 11943 32969
rect 11885 32929 11897 32963
rect 11931 32960 11943 32963
rect 12894 32960 12900 32972
rect 11931 32932 12900 32960
rect 11931 32929 11943 32932
rect 11885 32923 11943 32929
rect 12894 32920 12900 32932
rect 12952 32920 12958 32972
rect 15120 32960 15148 33000
rect 15562 32988 15568 33000
rect 15620 32988 15626 33040
rect 15028 32932 15148 32960
rect 9732 32864 10272 32892
rect 10965 32895 11023 32901
rect 9732 32852 9738 32864
rect 10965 32861 10977 32895
rect 11011 32892 11023 32895
rect 11238 32892 11244 32904
rect 11011 32864 11244 32892
rect 11011 32861 11023 32864
rect 10965 32855 11023 32861
rect 11238 32852 11244 32864
rect 11296 32892 11302 32904
rect 12342 32892 12348 32904
rect 11296 32864 12348 32892
rect 11296 32852 11302 32864
rect 12342 32852 12348 32864
rect 12400 32852 12406 32904
rect 12434 32852 12440 32904
rect 12492 32892 12498 32904
rect 15028 32901 15056 32932
rect 15194 32920 15200 32972
rect 15252 32960 15258 32972
rect 15841 32963 15899 32969
rect 15252 32932 15297 32960
rect 15252 32920 15258 32932
rect 15841 32929 15853 32963
rect 15887 32960 15899 32963
rect 16666 32960 16672 32972
rect 15887 32932 16672 32960
rect 15887 32929 15899 32932
rect 15841 32923 15899 32929
rect 16666 32920 16672 32932
rect 16724 32920 16730 32972
rect 18414 32920 18420 32972
rect 18472 32960 18478 32972
rect 18708 32969 18736 33068
rect 19518 33056 19524 33068
rect 19576 33056 19582 33108
rect 19794 33056 19800 33108
rect 19852 33096 19858 33108
rect 19852 33068 21220 33096
rect 19852 33056 19858 33068
rect 21192 33037 21220 33068
rect 24210 33056 24216 33108
rect 24268 33096 24274 33108
rect 24581 33099 24639 33105
rect 24581 33096 24593 33099
rect 24268 33068 24593 33096
rect 24268 33056 24274 33068
rect 24581 33065 24593 33068
rect 24627 33065 24639 33099
rect 24581 33059 24639 33065
rect 26053 33099 26111 33105
rect 26053 33065 26065 33099
rect 26099 33096 26111 33099
rect 26234 33096 26240 33108
rect 26099 33068 26240 33096
rect 26099 33065 26111 33068
rect 26053 33059 26111 33065
rect 26234 33056 26240 33068
rect 26292 33056 26298 33108
rect 26602 33056 26608 33108
rect 26660 33096 26666 33108
rect 26697 33099 26755 33105
rect 26697 33096 26709 33099
rect 26660 33068 26709 33096
rect 26660 33056 26666 33068
rect 26697 33065 26709 33068
rect 26743 33065 26755 33099
rect 30098 33096 30104 33108
rect 26697 33059 26755 33065
rect 27724 33068 30104 33096
rect 27724 33040 27752 33068
rect 30098 33056 30104 33068
rect 30156 33056 30162 33108
rect 30374 33056 30380 33108
rect 30432 33096 30438 33108
rect 30469 33099 30527 33105
rect 30469 33096 30481 33099
rect 30432 33068 30481 33096
rect 30432 33056 30438 33068
rect 30469 33065 30481 33068
rect 30515 33065 30527 33099
rect 30469 33059 30527 33065
rect 34333 33099 34391 33105
rect 34333 33065 34345 33099
rect 34379 33096 34391 33099
rect 34514 33096 34520 33108
rect 34379 33068 34520 33096
rect 34379 33065 34391 33068
rect 34333 33059 34391 33065
rect 34514 33056 34520 33068
rect 34572 33056 34578 33108
rect 21177 33031 21235 33037
rect 21177 32997 21189 33031
rect 21223 33028 21235 33031
rect 27706 33028 27712 33040
rect 21223 33000 27568 33028
rect 27667 33000 27712 33028
rect 21223 32997 21235 33000
rect 21177 32991 21235 32997
rect 18601 32963 18659 32969
rect 18601 32960 18613 32963
rect 18472 32932 18613 32960
rect 18472 32920 18478 32932
rect 18601 32929 18613 32932
rect 18647 32929 18659 32963
rect 18601 32923 18659 32929
rect 18693 32963 18751 32969
rect 18693 32929 18705 32963
rect 18739 32929 18751 32963
rect 18693 32923 18751 32929
rect 19429 32963 19487 32969
rect 19429 32929 19441 32963
rect 19475 32960 19487 32963
rect 22094 32960 22100 32972
rect 19475 32932 22100 32960
rect 19475 32929 19487 32932
rect 19429 32923 19487 32929
rect 13265 32895 13323 32901
rect 13265 32892 13277 32895
rect 12492 32864 13277 32892
rect 12492 32852 12498 32864
rect 13265 32861 13277 32864
rect 13311 32861 13323 32895
rect 13265 32855 13323 32861
rect 15013 32895 15071 32901
rect 15013 32861 15025 32895
rect 15059 32861 15071 32895
rect 15013 32855 15071 32861
rect 17954 32852 17960 32904
rect 18012 32892 18018 32904
rect 18708 32892 18736 32923
rect 22094 32920 22100 32932
rect 22152 32960 22158 32972
rect 22557 32963 22615 32969
rect 22557 32960 22569 32963
rect 22152 32932 22569 32960
rect 22152 32920 22158 32932
rect 22557 32929 22569 32932
rect 22603 32929 22615 32963
rect 22557 32923 22615 32929
rect 23753 32963 23811 32969
rect 23753 32929 23765 32963
rect 23799 32960 23811 32963
rect 23934 32960 23940 32972
rect 23799 32932 23940 32960
rect 23799 32929 23811 32932
rect 23753 32923 23811 32929
rect 23934 32920 23940 32932
rect 23992 32920 23998 32972
rect 25130 32960 25136 32972
rect 25091 32932 25136 32960
rect 25130 32920 25136 32932
rect 25188 32920 25194 32972
rect 26694 32920 26700 32972
rect 26752 32960 26758 32972
rect 27433 32963 27491 32969
rect 27433 32960 27445 32963
rect 26752 32932 27445 32960
rect 26752 32920 26758 32932
rect 27433 32929 27445 32932
rect 27479 32929 27491 32963
rect 27433 32923 27491 32929
rect 21818 32892 21824 32904
rect 18012 32864 18736 32892
rect 21779 32864 21824 32892
rect 18012 32852 18018 32864
rect 21818 32852 21824 32864
rect 21876 32852 21882 32904
rect 23569 32895 23627 32901
rect 23569 32861 23581 32895
rect 23615 32892 23627 32895
rect 23842 32892 23848 32904
rect 23615 32864 23848 32892
rect 23615 32861 23627 32864
rect 23569 32855 23627 32861
rect 23842 32852 23848 32864
rect 23900 32892 23906 32904
rect 25041 32895 25099 32901
rect 25041 32892 25053 32895
rect 23900 32864 25053 32892
rect 23900 32852 23906 32864
rect 25041 32861 25053 32864
rect 25087 32861 25099 32895
rect 25041 32855 25099 32861
rect 26145 32895 26203 32901
rect 26145 32861 26157 32895
rect 26191 32892 26203 32895
rect 26602 32892 26608 32904
rect 26191 32864 26608 32892
rect 26191 32861 26203 32864
rect 26145 32855 26203 32861
rect 26602 32852 26608 32864
rect 26660 32892 26666 32904
rect 26789 32895 26847 32901
rect 26789 32892 26801 32895
rect 26660 32864 26801 32892
rect 26660 32852 26666 32864
rect 26789 32861 26801 32864
rect 26835 32861 26847 32895
rect 26789 32855 26847 32861
rect 7282 32784 7288 32836
rect 7340 32824 7346 32836
rect 9953 32827 10011 32833
rect 7340 32796 7498 32824
rect 7340 32784 7346 32796
rect 9953 32793 9965 32827
rect 9999 32824 10011 32827
rect 12158 32824 12164 32836
rect 9999 32796 12164 32824
rect 9999 32793 10011 32796
rect 9953 32787 10011 32793
rect 12158 32784 12164 32796
rect 12216 32784 12222 32836
rect 16850 32784 16856 32836
rect 16908 32784 16914 32836
rect 18874 32784 18880 32836
rect 18932 32824 18938 32836
rect 19705 32827 19763 32833
rect 19705 32824 19717 32827
rect 18932 32796 19717 32824
rect 18932 32784 18938 32796
rect 19705 32793 19717 32796
rect 19751 32793 19763 32827
rect 19705 32787 19763 32793
rect 20438 32784 20444 32836
rect 20496 32784 20502 32836
rect 23661 32827 23719 32833
rect 23661 32793 23673 32827
rect 23707 32824 23719 32827
rect 25314 32824 25320 32836
rect 23707 32796 25320 32824
rect 23707 32793 23719 32796
rect 23661 32787 23719 32793
rect 25314 32784 25320 32796
rect 25372 32784 25378 32836
rect 27540 32824 27568 33000
rect 27706 32988 27712 33000
rect 27764 32988 27770 33040
rect 27893 33031 27951 33037
rect 27893 32997 27905 33031
rect 27939 33028 27951 33031
rect 30006 33028 30012 33040
rect 27939 33000 30012 33028
rect 27939 32997 27951 33000
rect 27893 32991 27951 32997
rect 30006 32988 30012 33000
rect 30064 32988 30070 33040
rect 28350 32920 28356 32972
rect 28408 32960 28414 32972
rect 28445 32963 28503 32969
rect 28445 32960 28457 32963
rect 28408 32932 28457 32960
rect 28408 32920 28414 32932
rect 28445 32929 28457 32932
rect 28491 32929 28503 32963
rect 28445 32923 28503 32929
rect 28537 32963 28595 32969
rect 28537 32929 28549 32963
rect 28583 32960 28595 32963
rect 29178 32960 29184 32972
rect 28583 32932 29184 32960
rect 28583 32929 28595 32932
rect 28537 32923 28595 32929
rect 29178 32920 29184 32932
rect 29236 32920 29242 32972
rect 30116 32969 30144 33056
rect 31021 33031 31079 33037
rect 31021 32997 31033 33031
rect 31067 33028 31079 33031
rect 31294 33028 31300 33040
rect 31067 33000 31300 33028
rect 31067 32997 31079 33000
rect 31021 32991 31079 32997
rect 31294 32988 31300 33000
rect 31352 32988 31358 33040
rect 31386 32988 31392 33040
rect 31444 32988 31450 33040
rect 30101 32963 30159 32969
rect 30101 32929 30113 32963
rect 30147 32929 30159 32963
rect 31404 32960 31432 32988
rect 30101 32923 30159 32929
rect 30300 32932 31432 32960
rect 27982 32852 27988 32904
rect 28040 32892 28046 32904
rect 28626 32892 28632 32904
rect 28040 32864 28632 32892
rect 28040 32852 28046 32864
rect 28626 32852 28632 32864
rect 28684 32852 28690 32904
rect 28721 32895 28779 32901
rect 28721 32861 28733 32895
rect 28767 32892 28779 32895
rect 29362 32892 29368 32904
rect 28767 32864 29368 32892
rect 28767 32861 28779 32864
rect 28721 32855 28779 32861
rect 29362 32852 29368 32864
rect 29420 32852 29426 32904
rect 30300 32901 30328 32932
rect 33502 32920 33508 32972
rect 33560 32960 33566 32972
rect 33689 32963 33747 32969
rect 33689 32960 33701 32963
rect 33560 32932 33701 32960
rect 33560 32920 33566 32932
rect 33689 32929 33701 32932
rect 33735 32929 33747 32963
rect 33689 32923 33747 32929
rect 30285 32895 30343 32901
rect 30285 32861 30297 32895
rect 30331 32861 30343 32895
rect 30285 32855 30343 32861
rect 32766 32852 32772 32904
rect 32824 32892 32830 32904
rect 32824 32864 32869 32892
rect 32824 32852 32830 32864
rect 27540 32796 31156 32824
rect 11054 32756 11060 32768
rect 11015 32728 11060 32756
rect 11054 32716 11060 32728
rect 11112 32716 11118 32768
rect 11514 32716 11520 32768
rect 11572 32756 11578 32768
rect 11977 32759 12035 32765
rect 11977 32756 11989 32759
rect 11572 32728 11989 32756
rect 11572 32716 11578 32728
rect 11977 32725 11989 32728
rect 12023 32725 12035 32759
rect 11977 32719 12035 32725
rect 13173 32759 13231 32765
rect 13173 32725 13185 32759
rect 13219 32756 13231 32759
rect 13354 32756 13360 32768
rect 13219 32728 13360 32756
rect 13219 32725 13231 32728
rect 13173 32719 13231 32725
rect 13354 32716 13360 32728
rect 13412 32716 13418 32768
rect 15105 32759 15163 32765
rect 15105 32725 15117 32759
rect 15151 32756 15163 32759
rect 15194 32756 15200 32768
rect 15151 32728 15200 32756
rect 15151 32725 15163 32728
rect 15105 32719 15163 32725
rect 15194 32716 15200 32728
rect 15252 32756 15258 32768
rect 16022 32756 16028 32768
rect 15252 32728 16028 32756
rect 15252 32716 15258 32728
rect 16022 32716 16028 32728
rect 16080 32716 16086 32768
rect 17494 32716 17500 32768
rect 17552 32756 17558 32768
rect 17589 32759 17647 32765
rect 17589 32756 17601 32759
rect 17552 32728 17601 32756
rect 17552 32716 17558 32728
rect 17589 32725 17601 32728
rect 17635 32756 17647 32759
rect 17862 32756 17868 32768
rect 17635 32728 17868 32756
rect 17635 32725 17647 32728
rect 17589 32719 17647 32725
rect 17862 32716 17868 32728
rect 17920 32716 17926 32768
rect 18506 32756 18512 32768
rect 18467 32728 18512 32756
rect 18506 32716 18512 32728
rect 18564 32716 18570 32768
rect 23198 32756 23204 32768
rect 23159 32728 23204 32756
rect 23198 32716 23204 32728
rect 23256 32716 23262 32768
rect 24946 32756 24952 32768
rect 24907 32728 24952 32756
rect 24946 32716 24952 32728
rect 25004 32716 25010 32768
rect 28258 32716 28264 32768
rect 28316 32756 28322 32768
rect 28905 32759 28963 32765
rect 28905 32756 28917 32759
rect 28316 32728 28917 32756
rect 28316 32716 28322 32728
rect 28905 32725 28917 32728
rect 28951 32725 28963 32759
rect 31128 32756 31156 32796
rect 32030 32784 32036 32836
rect 32088 32784 32094 32836
rect 32493 32827 32551 32833
rect 32493 32793 32505 32827
rect 32539 32824 32551 32827
rect 33042 32824 33048 32836
rect 32539 32796 33048 32824
rect 32539 32793 32551 32796
rect 32493 32787 32551 32793
rect 33042 32784 33048 32796
rect 33100 32784 33106 32836
rect 33134 32784 33140 32836
rect 33192 32824 33198 32836
rect 33965 32827 34023 32833
rect 33965 32824 33977 32827
rect 33192 32796 33977 32824
rect 33192 32784 33198 32796
rect 33965 32793 33977 32796
rect 34011 32793 34023 32827
rect 33965 32787 34023 32793
rect 33873 32759 33931 32765
rect 33873 32756 33885 32759
rect 31128 32728 33885 32756
rect 28905 32719 28963 32725
rect 33873 32725 33885 32728
rect 33919 32725 33931 32759
rect 33873 32719 33931 32725
rect 1104 32666 37628 32688
rect 1104 32614 4874 32666
rect 4926 32614 4938 32666
rect 4990 32614 5002 32666
rect 5054 32614 5066 32666
rect 5118 32614 5130 32666
rect 5182 32614 35594 32666
rect 35646 32614 35658 32666
rect 35710 32614 35722 32666
rect 35774 32614 35786 32666
rect 35838 32614 35850 32666
rect 35902 32614 37628 32666
rect 1104 32592 37628 32614
rect 7377 32555 7435 32561
rect 7377 32521 7389 32555
rect 7423 32552 7435 32555
rect 8110 32552 8116 32564
rect 7423 32524 8116 32552
rect 7423 32521 7435 32524
rect 7377 32515 7435 32521
rect 8110 32512 8116 32524
rect 8168 32512 8174 32564
rect 9398 32552 9404 32564
rect 8404 32524 9404 32552
rect 7929 32487 7987 32493
rect 7929 32453 7941 32487
rect 7975 32484 7987 32487
rect 8294 32484 8300 32496
rect 7975 32456 8300 32484
rect 7975 32453 7987 32456
rect 7929 32447 7987 32453
rect 8294 32444 8300 32456
rect 8352 32444 8358 32496
rect 6549 32419 6607 32425
rect 6549 32385 6561 32419
rect 6595 32416 6607 32419
rect 7193 32419 7251 32425
rect 6595 32388 6914 32416
rect 6595 32385 6607 32388
rect 6549 32379 6607 32385
rect 6886 32348 6914 32388
rect 7193 32385 7205 32419
rect 7239 32416 7251 32419
rect 8021 32419 8079 32425
rect 7239 32388 7972 32416
rect 7239 32385 7251 32388
rect 7193 32379 7251 32385
rect 7834 32348 7840 32360
rect 6886 32320 7840 32348
rect 7834 32308 7840 32320
rect 7892 32308 7898 32360
rect 7944 32348 7972 32388
rect 8021 32385 8033 32419
rect 8067 32416 8079 32419
rect 8404 32416 8432 32524
rect 9398 32512 9404 32524
rect 9456 32512 9462 32564
rect 14093 32555 14151 32561
rect 14093 32521 14105 32555
rect 14139 32552 14151 32555
rect 15194 32552 15200 32564
rect 14139 32524 15200 32552
rect 14139 32521 14151 32524
rect 14093 32515 14151 32521
rect 15194 32512 15200 32524
rect 15252 32512 15258 32564
rect 18506 32512 18512 32564
rect 18564 32552 18570 32564
rect 19153 32555 19211 32561
rect 19153 32552 19165 32555
rect 18564 32524 19165 32552
rect 18564 32512 18570 32524
rect 19153 32521 19165 32524
rect 19199 32521 19211 32555
rect 19153 32515 19211 32521
rect 19613 32555 19671 32561
rect 19613 32521 19625 32555
rect 19659 32552 19671 32555
rect 19794 32552 19800 32564
rect 19659 32524 19800 32552
rect 19659 32521 19671 32524
rect 19613 32515 19671 32521
rect 19794 32512 19800 32524
rect 19852 32512 19858 32564
rect 20438 32552 20444 32564
rect 20399 32524 20444 32552
rect 20438 32512 20444 32524
rect 20496 32512 20502 32564
rect 22278 32512 22284 32564
rect 22336 32552 22342 32564
rect 22649 32555 22707 32561
rect 22649 32552 22661 32555
rect 22336 32524 22661 32552
rect 22336 32512 22342 32524
rect 22649 32521 22661 32524
rect 22695 32521 22707 32555
rect 22649 32515 22707 32521
rect 23382 32512 23388 32564
rect 23440 32552 23446 32564
rect 23661 32555 23719 32561
rect 23661 32552 23673 32555
rect 23440 32524 23673 32552
rect 23440 32512 23446 32524
rect 23661 32521 23673 32524
rect 23707 32552 23719 32555
rect 24765 32555 24823 32561
rect 24765 32552 24777 32555
rect 23707 32524 24777 32552
rect 23707 32521 23719 32524
rect 23661 32515 23719 32521
rect 24765 32521 24777 32524
rect 24811 32521 24823 32555
rect 24765 32515 24823 32521
rect 25225 32555 25283 32561
rect 25225 32521 25237 32555
rect 25271 32521 25283 32555
rect 25225 32515 25283 32521
rect 11054 32444 11060 32496
rect 11112 32484 11118 32496
rect 25130 32484 25136 32496
rect 11112 32456 14398 32484
rect 24688 32456 25136 32484
rect 11112 32444 11118 32456
rect 8067 32388 8432 32416
rect 8481 32419 8539 32425
rect 8067 32385 8079 32388
rect 8021 32379 8079 32385
rect 8481 32385 8493 32419
rect 8527 32416 8539 32419
rect 8938 32416 8944 32428
rect 8527 32388 8944 32416
rect 8527 32385 8539 32388
rect 8481 32379 8539 32385
rect 8938 32376 8944 32388
rect 8996 32376 9002 32428
rect 9306 32416 9312 32428
rect 9267 32388 9312 32416
rect 9306 32376 9312 32388
rect 9364 32416 9370 32428
rect 10321 32419 10379 32425
rect 10321 32416 10333 32419
rect 9364 32388 10333 32416
rect 9364 32376 9370 32388
rect 10321 32385 10333 32388
rect 10367 32385 10379 32419
rect 10962 32416 10968 32428
rect 10923 32388 10968 32416
rect 10321 32379 10379 32385
rect 10962 32376 10968 32388
rect 11020 32376 11026 32428
rect 12066 32416 12072 32428
rect 12027 32388 12072 32416
rect 12066 32376 12072 32388
rect 12124 32376 12130 32428
rect 12342 32376 12348 32428
rect 12400 32416 12406 32428
rect 13357 32419 13415 32425
rect 13357 32416 13369 32419
rect 12400 32388 13369 32416
rect 12400 32376 12406 32388
rect 13357 32385 13369 32388
rect 13403 32385 13415 32419
rect 13357 32379 13415 32385
rect 16850 32376 16856 32428
rect 16908 32416 16914 32428
rect 17037 32419 17095 32425
rect 17037 32416 17049 32419
rect 16908 32388 17049 32416
rect 16908 32376 16914 32388
rect 17037 32385 17049 32388
rect 17083 32385 17095 32419
rect 18046 32416 18052 32428
rect 18007 32388 18052 32416
rect 17037 32379 17095 32385
rect 18046 32376 18052 32388
rect 18104 32376 18110 32428
rect 19518 32416 19524 32428
rect 19479 32388 19524 32416
rect 19518 32376 19524 32388
rect 19576 32376 19582 32428
rect 20349 32419 20407 32425
rect 20349 32385 20361 32419
rect 20395 32385 20407 32419
rect 21266 32416 21272 32428
rect 21227 32388 21272 32416
rect 20349 32379 20407 32385
rect 9122 32348 9128 32360
rect 7944 32320 9128 32348
rect 9122 32308 9128 32320
rect 9180 32308 9186 32360
rect 12158 32348 12164 32360
rect 12119 32320 12164 32348
rect 12158 32308 12164 32320
rect 12216 32308 12222 32360
rect 12253 32351 12311 32357
rect 12253 32317 12265 32351
rect 12299 32348 12311 32351
rect 12618 32348 12624 32360
rect 12299 32320 12624 32348
rect 12299 32317 12311 32320
rect 12253 32311 12311 32317
rect 12618 32308 12624 32320
rect 12676 32308 12682 32360
rect 13449 32351 13507 32357
rect 13449 32317 13461 32351
rect 13495 32348 13507 32351
rect 15194 32348 15200 32360
rect 13495 32320 15200 32348
rect 13495 32317 13507 32320
rect 13449 32311 13507 32317
rect 15194 32308 15200 32320
rect 15252 32308 15258 32360
rect 15841 32351 15899 32357
rect 15841 32317 15853 32351
rect 15887 32348 15899 32351
rect 16666 32348 16672 32360
rect 15887 32320 16672 32348
rect 15887 32317 15899 32320
rect 15841 32311 15899 32317
rect 16666 32308 16672 32320
rect 16724 32348 16730 32360
rect 17126 32348 17132 32360
rect 16724 32320 17132 32348
rect 16724 32308 16730 32320
rect 17126 32308 17132 32320
rect 17184 32308 17190 32360
rect 19702 32308 19708 32360
rect 19760 32348 19766 32360
rect 19760 32320 19805 32348
rect 19760 32308 19766 32320
rect 20070 32308 20076 32360
rect 20128 32348 20134 32360
rect 20364 32348 20392 32379
rect 21266 32376 21272 32388
rect 21324 32376 21330 32428
rect 22186 32416 22192 32428
rect 22147 32388 22192 32416
rect 22186 32376 22192 32388
rect 22244 32376 22250 32428
rect 22830 32416 22836 32428
rect 22791 32388 22836 32416
rect 22830 32376 22836 32388
rect 22888 32376 22894 32428
rect 20898 32348 20904 32360
rect 20128 32320 20904 32348
rect 20128 32308 20134 32320
rect 20898 32308 20904 32320
rect 20956 32348 20962 32360
rect 22278 32348 22284 32360
rect 20956 32320 22284 32348
rect 20956 32308 20962 32320
rect 22278 32308 22284 32320
rect 22336 32308 22342 32360
rect 23753 32351 23811 32357
rect 23753 32317 23765 32351
rect 23799 32317 23811 32351
rect 23934 32348 23940 32360
rect 23895 32320 23940 32348
rect 23753 32311 23811 32317
rect 12176 32280 12204 32308
rect 12342 32280 12348 32292
rect 12176 32252 12348 32280
rect 12342 32240 12348 32252
rect 12400 32240 12406 32292
rect 23768 32280 23796 32311
rect 23934 32308 23940 32320
rect 23992 32308 23998 32360
rect 24688 32357 24716 32456
rect 25130 32444 25136 32456
rect 25188 32444 25194 32496
rect 24857 32419 24915 32425
rect 24857 32385 24869 32419
rect 24903 32385 24915 32419
rect 25240 32416 25268 32515
rect 28994 32512 29000 32564
rect 29052 32552 29058 32564
rect 29546 32552 29552 32564
rect 29052 32524 29552 32552
rect 29052 32512 29058 32524
rect 29546 32512 29552 32524
rect 29604 32552 29610 32564
rect 30101 32555 30159 32561
rect 30101 32552 30113 32555
rect 29604 32524 30113 32552
rect 29604 32512 29610 32524
rect 30101 32521 30113 32524
rect 30147 32521 30159 32555
rect 30101 32515 30159 32521
rect 30926 32512 30932 32564
rect 30984 32552 30990 32564
rect 31205 32555 31263 32561
rect 31205 32552 31217 32555
rect 30984 32524 31217 32552
rect 30984 32512 30990 32524
rect 31205 32521 31217 32524
rect 31251 32521 31263 32555
rect 33042 32552 33048 32564
rect 33003 32524 33048 32552
rect 31205 32515 31263 32521
rect 33042 32512 33048 32524
rect 33100 32512 33106 32564
rect 27522 32444 27528 32496
rect 27580 32484 27586 32496
rect 27801 32487 27859 32493
rect 27801 32484 27813 32487
rect 27580 32456 27813 32484
rect 27580 32444 27586 32456
rect 27801 32453 27813 32456
rect 27847 32453 27859 32487
rect 29638 32484 29644 32496
rect 29599 32456 29644 32484
rect 27801 32447 27859 32453
rect 25869 32419 25927 32425
rect 25869 32416 25881 32419
rect 25240 32388 25881 32416
rect 24857 32379 24915 32385
rect 25869 32385 25881 32388
rect 25915 32385 25927 32419
rect 25869 32379 25927 32385
rect 26513 32419 26571 32425
rect 26513 32385 26525 32419
rect 26559 32416 26571 32419
rect 26602 32416 26608 32428
rect 26559 32388 26608 32416
rect 26559 32385 26571 32388
rect 26513 32379 26571 32385
rect 24673 32351 24731 32357
rect 24673 32317 24685 32351
rect 24719 32317 24731 32351
rect 24872 32348 24900 32379
rect 26602 32376 26608 32388
rect 26660 32376 26666 32428
rect 27341 32419 27399 32425
rect 27341 32385 27353 32419
rect 27387 32416 27399 32419
rect 27706 32416 27712 32428
rect 27387 32388 27712 32416
rect 27387 32385 27399 32388
rect 27341 32379 27399 32385
rect 27706 32376 27712 32388
rect 27764 32376 27770 32428
rect 25314 32348 25320 32360
rect 24872 32320 25320 32348
rect 24673 32311 24731 32317
rect 25314 32308 25320 32320
rect 25372 32308 25378 32360
rect 25038 32280 25044 32292
rect 23768 32252 25044 32280
rect 25038 32240 25044 32252
rect 25096 32240 25102 32292
rect 6638 32172 6644 32224
rect 6696 32212 6702 32224
rect 6733 32215 6791 32221
rect 6733 32212 6745 32215
rect 6696 32184 6745 32212
rect 6696 32172 6702 32184
rect 6733 32181 6745 32184
rect 6779 32181 6791 32215
rect 8662 32212 8668 32224
rect 8623 32184 8668 32212
rect 6733 32175 6791 32181
rect 8662 32172 8668 32184
rect 8720 32172 8726 32224
rect 9214 32212 9220 32224
rect 9175 32184 9220 32212
rect 9214 32172 9220 32184
rect 9272 32172 9278 32224
rect 10413 32215 10471 32221
rect 10413 32181 10425 32215
rect 10459 32212 10471 32215
rect 10502 32212 10508 32224
rect 10459 32184 10508 32212
rect 10459 32181 10471 32184
rect 10413 32175 10471 32181
rect 10502 32172 10508 32184
rect 10560 32172 10566 32224
rect 11146 32212 11152 32224
rect 11107 32184 11152 32212
rect 11146 32172 11152 32184
rect 11204 32172 11210 32224
rect 11698 32212 11704 32224
rect 11659 32184 11704 32212
rect 11698 32172 11704 32184
rect 11756 32172 11762 32224
rect 14458 32172 14464 32224
rect 14516 32212 14522 32224
rect 15577 32215 15635 32221
rect 15577 32212 15589 32215
rect 14516 32184 15589 32212
rect 14516 32172 14522 32184
rect 15577 32181 15589 32184
rect 15623 32181 15635 32215
rect 15577 32175 15635 32181
rect 16853 32215 16911 32221
rect 16853 32181 16865 32215
rect 16899 32212 16911 32215
rect 17310 32212 17316 32224
rect 16899 32184 17316 32212
rect 16899 32181 16911 32184
rect 16853 32175 16911 32181
rect 17310 32172 17316 32184
rect 17368 32172 17374 32224
rect 18141 32215 18199 32221
rect 18141 32181 18153 32215
rect 18187 32212 18199 32215
rect 18506 32212 18512 32224
rect 18187 32184 18512 32212
rect 18187 32181 18199 32184
rect 18141 32175 18199 32181
rect 18506 32172 18512 32184
rect 18564 32172 18570 32224
rect 21361 32215 21419 32221
rect 21361 32181 21373 32215
rect 21407 32212 21419 32215
rect 21450 32212 21456 32224
rect 21407 32184 21456 32212
rect 21407 32181 21419 32184
rect 21361 32175 21419 32181
rect 21450 32172 21456 32184
rect 21508 32172 21514 32224
rect 22002 32212 22008 32224
rect 21963 32184 22008 32212
rect 22002 32172 22008 32184
rect 22060 32172 22066 32224
rect 23290 32212 23296 32224
rect 23251 32184 23296 32212
rect 23290 32172 23296 32184
rect 23348 32172 23354 32224
rect 24946 32172 24952 32224
rect 25004 32212 25010 32224
rect 25685 32215 25743 32221
rect 25685 32212 25697 32215
rect 25004 32184 25697 32212
rect 25004 32172 25010 32184
rect 25685 32181 25697 32184
rect 25731 32181 25743 32215
rect 26418 32212 26424 32224
rect 26379 32184 26424 32212
rect 25685 32175 25743 32181
rect 26418 32172 26424 32184
rect 26476 32172 26482 32224
rect 27249 32215 27307 32221
rect 27249 32181 27261 32215
rect 27295 32212 27307 32215
rect 27706 32212 27712 32224
rect 27295 32184 27712 32212
rect 27295 32181 27307 32184
rect 27249 32175 27307 32181
rect 27706 32172 27712 32184
rect 27764 32172 27770 32224
rect 27816 32212 27844 32447
rect 29638 32444 29644 32456
rect 29696 32444 29702 32496
rect 31128 32456 31754 32484
rect 31128 32428 31156 32456
rect 29914 32416 29920 32428
rect 28276 32388 29920 32416
rect 28276 32357 28304 32388
rect 29914 32376 29920 32388
rect 29972 32376 29978 32428
rect 31110 32416 31116 32428
rect 31071 32388 31116 32416
rect 31110 32376 31116 32388
rect 31168 32376 31174 32428
rect 31294 32376 31300 32428
rect 31352 32416 31358 32428
rect 31389 32419 31447 32425
rect 31389 32416 31401 32419
rect 31352 32388 31401 32416
rect 31352 32376 31358 32388
rect 31389 32385 31401 32388
rect 31435 32385 31447 32419
rect 31726 32416 31754 32456
rect 32030 32444 32036 32496
rect 32088 32484 32094 32496
rect 34333 32487 34391 32493
rect 34333 32484 34345 32487
rect 32088 32456 34345 32484
rect 32088 32444 32094 32456
rect 34333 32453 34345 32456
rect 34379 32453 34391 32487
rect 34333 32447 34391 32453
rect 32493 32419 32551 32425
rect 32493 32416 32505 32419
rect 31726 32388 32505 32416
rect 31389 32379 31447 32385
rect 32493 32385 32505 32388
rect 32539 32385 32551 32419
rect 32493 32379 32551 32385
rect 32953 32419 33011 32425
rect 32953 32385 32965 32419
rect 32999 32385 33011 32419
rect 32953 32379 33011 32385
rect 33137 32419 33195 32425
rect 33137 32385 33149 32419
rect 33183 32385 33195 32419
rect 33778 32416 33784 32428
rect 33739 32388 33784 32416
rect 33137 32379 33195 32385
rect 28261 32351 28319 32357
rect 28261 32317 28273 32351
rect 28307 32317 28319 32351
rect 28261 32311 28319 32317
rect 28721 32351 28779 32357
rect 28721 32317 28733 32351
rect 28767 32348 28779 32351
rect 29181 32351 29239 32357
rect 28767 32320 29132 32348
rect 28767 32317 28779 32320
rect 28721 32311 28779 32317
rect 28169 32283 28227 32289
rect 28169 32249 28181 32283
rect 28215 32280 28227 32283
rect 28736 32280 28764 32311
rect 28215 32252 28764 32280
rect 28997 32283 29055 32289
rect 28215 32249 28227 32252
rect 28169 32243 28227 32249
rect 28997 32249 29009 32283
rect 29043 32249 29055 32283
rect 29104 32280 29132 32320
rect 29181 32317 29193 32351
rect 29227 32348 29239 32351
rect 29733 32351 29791 32357
rect 29733 32348 29745 32351
rect 29227 32320 29745 32348
rect 29227 32317 29239 32320
rect 29181 32311 29239 32317
rect 29733 32317 29745 32320
rect 29779 32317 29791 32351
rect 32968 32348 32996 32379
rect 29733 32311 29791 32317
rect 31726 32320 32996 32348
rect 31294 32280 31300 32292
rect 29104 32252 31300 32280
rect 28997 32243 29055 32249
rect 29012 32212 29040 32243
rect 31294 32240 31300 32252
rect 31352 32240 31358 32292
rect 31389 32283 31447 32289
rect 31389 32249 31401 32283
rect 31435 32280 31447 32283
rect 31726 32280 31754 32320
rect 32398 32280 32404 32292
rect 31435 32252 31754 32280
rect 32359 32252 32404 32280
rect 31435 32249 31447 32252
rect 31389 32243 31447 32249
rect 32398 32240 32404 32252
rect 32456 32240 32462 32292
rect 27816 32184 29040 32212
rect 29917 32215 29975 32221
rect 29917 32181 29929 32215
rect 29963 32212 29975 32215
rect 30006 32212 30012 32224
rect 29963 32184 30012 32212
rect 29963 32181 29975 32184
rect 29917 32175 29975 32181
rect 30006 32172 30012 32184
rect 30064 32172 30070 32224
rect 30834 32172 30840 32224
rect 30892 32212 30898 32224
rect 31478 32212 31484 32224
rect 30892 32184 31484 32212
rect 30892 32172 30898 32184
rect 31478 32172 31484 32184
rect 31536 32212 31542 32224
rect 33152 32212 33180 32379
rect 33778 32376 33784 32388
rect 33836 32416 33842 32428
rect 34241 32419 34299 32425
rect 34241 32416 34253 32419
rect 33836 32388 34253 32416
rect 33836 32376 33842 32388
rect 34241 32385 34253 32388
rect 34287 32385 34299 32419
rect 34241 32379 34299 32385
rect 33686 32212 33692 32224
rect 31536 32184 33180 32212
rect 33647 32184 33692 32212
rect 31536 32172 31542 32184
rect 33686 32172 33692 32184
rect 33744 32172 33750 32224
rect 1104 32122 37628 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 37628 32122
rect 1104 32048 37628 32070
rect 7282 32008 7288 32020
rect 7243 31980 7288 32008
rect 7282 31968 7288 31980
rect 7340 31968 7346 32020
rect 7834 32008 7840 32020
rect 7795 31980 7840 32008
rect 7834 31968 7840 31980
rect 7892 31968 7898 32020
rect 9309 32011 9367 32017
rect 9309 31977 9321 32011
rect 9355 32008 9367 32011
rect 11054 32008 11060 32020
rect 9355 31980 11060 32008
rect 9355 31977 9367 31980
rect 9309 31971 9367 31977
rect 11054 31968 11060 31980
rect 11112 31968 11118 32020
rect 11146 31968 11152 32020
rect 11204 32008 11210 32020
rect 12234 32011 12292 32017
rect 12234 32008 12246 32011
rect 11204 31980 12246 32008
rect 11204 31968 11210 31980
rect 12234 31977 12246 31980
rect 12280 31977 12292 32011
rect 12234 31971 12292 31977
rect 12342 31968 12348 32020
rect 12400 32008 12406 32020
rect 13725 32011 13783 32017
rect 13725 32008 13737 32011
rect 12400 31980 13737 32008
rect 12400 31968 12406 31980
rect 13725 31977 13737 31980
rect 13771 31977 13783 32011
rect 15010 32008 15016 32020
rect 14971 31980 15016 32008
rect 13725 31971 13783 31977
rect 11514 31940 11520 31952
rect 11475 31912 11520 31940
rect 11514 31900 11520 31912
rect 11572 31900 11578 31952
rect 13740 31940 13768 31971
rect 15010 31968 15016 31980
rect 15068 31968 15074 32020
rect 20980 32011 21038 32017
rect 20980 31977 20992 32011
rect 21026 32008 21038 32011
rect 22002 32008 22008 32020
rect 21026 31980 22008 32008
rect 21026 31977 21038 31980
rect 20980 31971 21038 31977
rect 22002 31968 22008 31980
rect 22060 31968 22066 32020
rect 22186 31968 22192 32020
rect 22244 32008 22250 32020
rect 22925 32011 22983 32017
rect 22925 32008 22937 32011
rect 22244 31980 22937 32008
rect 22244 31968 22250 31980
rect 22925 31977 22937 31980
rect 22971 31977 22983 32011
rect 22925 31971 22983 31977
rect 27801 32011 27859 32017
rect 27801 31977 27813 32011
rect 27847 32008 27859 32011
rect 29270 32008 29276 32020
rect 27847 31980 29276 32008
rect 27847 31977 27859 31980
rect 27801 31971 27859 31977
rect 29270 31968 29276 31980
rect 29328 31968 29334 32020
rect 30926 31968 30932 32020
rect 30984 32008 30990 32020
rect 33045 32011 33103 32017
rect 33045 32008 33057 32011
rect 30984 31980 33057 32008
rect 30984 31968 30990 31980
rect 33045 31977 33057 31980
rect 33091 31977 33103 32011
rect 33045 31971 33103 31977
rect 22094 31940 22100 31952
rect 13740 31912 14596 31940
rect 8018 31832 8024 31884
rect 8076 31872 8082 31884
rect 8389 31875 8447 31881
rect 8389 31872 8401 31875
rect 8076 31844 8401 31872
rect 8076 31832 8082 31844
rect 8389 31841 8401 31844
rect 8435 31841 8447 31875
rect 8389 31835 8447 31841
rect 8662 31832 8668 31884
rect 8720 31872 8726 31884
rect 10045 31875 10103 31881
rect 10045 31872 10057 31875
rect 8720 31844 10057 31872
rect 8720 31832 8726 31844
rect 10045 31841 10057 31844
rect 10091 31841 10103 31875
rect 10045 31835 10103 31841
rect 11977 31875 12035 31881
rect 11977 31841 11989 31875
rect 12023 31872 12035 31875
rect 12250 31872 12256 31884
rect 12023 31844 12256 31872
rect 12023 31841 12035 31844
rect 11977 31835 12035 31841
rect 12250 31832 12256 31844
rect 12308 31832 12314 31884
rect 14274 31832 14280 31884
rect 14332 31872 14338 31884
rect 14568 31881 14596 31912
rect 22066 31900 22100 31940
rect 22152 31900 22158 31952
rect 22465 31943 22523 31949
rect 22465 31909 22477 31943
rect 22511 31940 22523 31943
rect 23382 31940 23388 31952
rect 22511 31912 23388 31940
rect 22511 31909 22523 31912
rect 22465 31903 22523 31909
rect 23382 31900 23388 31912
rect 23440 31900 23446 31952
rect 29086 31940 29092 31952
rect 28736 31912 29092 31940
rect 14369 31875 14427 31881
rect 14369 31872 14381 31875
rect 14332 31844 14381 31872
rect 14332 31832 14338 31844
rect 14369 31841 14381 31844
rect 14415 31841 14427 31875
rect 14369 31835 14427 31841
rect 14553 31875 14611 31881
rect 14553 31841 14565 31875
rect 14599 31841 14611 31875
rect 16114 31872 16120 31884
rect 16075 31844 16120 31872
rect 14553 31835 14611 31841
rect 16114 31832 16120 31844
rect 16172 31832 16178 31884
rect 18877 31875 18935 31881
rect 18877 31841 18889 31875
rect 18923 31872 18935 31875
rect 19518 31872 19524 31884
rect 18923 31844 19524 31872
rect 18923 31841 18935 31844
rect 18877 31835 18935 31841
rect 19518 31832 19524 31844
rect 19576 31872 19582 31884
rect 19886 31872 19892 31884
rect 19576 31844 19892 31872
rect 19576 31832 19582 31844
rect 19886 31832 19892 31844
rect 19944 31832 19950 31884
rect 20717 31875 20775 31881
rect 20717 31841 20729 31875
rect 20763 31872 20775 31875
rect 22066 31872 22094 31900
rect 20763 31844 22094 31872
rect 20763 31841 20775 31844
rect 20717 31835 20775 31841
rect 22554 31832 22560 31884
rect 22612 31872 22618 31884
rect 23477 31875 23535 31881
rect 23477 31872 23489 31875
rect 22612 31844 23489 31872
rect 22612 31832 22618 31844
rect 23477 31841 23489 31844
rect 23523 31841 23535 31875
rect 24946 31872 24952 31884
rect 24907 31844 24952 31872
rect 23477 31835 23535 31841
rect 24946 31832 24952 31844
rect 25004 31832 25010 31884
rect 25314 31832 25320 31884
rect 25372 31872 25378 31884
rect 26421 31875 26479 31881
rect 26421 31872 26433 31875
rect 25372 31844 26433 31872
rect 25372 31832 25378 31844
rect 26421 31841 26433 31844
rect 26467 31872 26479 31875
rect 27890 31872 27896 31884
rect 26467 31844 27896 31872
rect 26467 31841 26479 31844
rect 26421 31835 26479 31841
rect 27890 31832 27896 31844
rect 27948 31832 27954 31884
rect 1765 31807 1823 31813
rect 1765 31773 1777 31807
rect 1811 31804 1823 31807
rect 1946 31804 1952 31816
rect 1811 31776 1952 31804
rect 1811 31773 1823 31776
rect 1765 31767 1823 31773
rect 1946 31764 1952 31776
rect 2004 31764 2010 31816
rect 6549 31807 6607 31813
rect 6549 31773 6561 31807
rect 6595 31804 6607 31807
rect 6914 31804 6920 31816
rect 6595 31776 6920 31804
rect 6595 31773 6607 31776
rect 6549 31767 6607 31773
rect 6914 31764 6920 31776
rect 6972 31804 6978 31816
rect 7098 31804 7104 31816
rect 6972 31776 7104 31804
rect 6972 31764 6978 31776
rect 7098 31764 7104 31776
rect 7156 31804 7162 31816
rect 7193 31807 7251 31813
rect 7193 31804 7205 31807
rect 7156 31776 7205 31804
rect 7156 31764 7162 31776
rect 7193 31773 7205 31776
rect 7239 31773 7251 31807
rect 9122 31804 9128 31816
rect 9083 31776 9128 31804
rect 7193 31767 7251 31773
rect 9122 31764 9128 31776
rect 9180 31764 9186 31816
rect 9766 31804 9772 31816
rect 9727 31776 9772 31804
rect 9766 31764 9772 31776
rect 9824 31764 9830 31816
rect 13354 31764 13360 31816
rect 13412 31764 13418 31816
rect 16022 31804 16028 31816
rect 15948 31776 16028 31804
rect 10502 31696 10508 31748
rect 10560 31696 10566 31748
rect 15948 31745 15976 31776
rect 16022 31764 16028 31776
rect 16080 31764 16086 31816
rect 17126 31804 17132 31816
rect 17039 31776 17132 31804
rect 17126 31764 17132 31776
rect 17184 31764 17190 31816
rect 18506 31764 18512 31816
rect 18564 31764 18570 31816
rect 19610 31804 19616 31816
rect 19571 31776 19616 31804
rect 19610 31764 19616 31776
rect 19668 31764 19674 31816
rect 20070 31804 20076 31816
rect 20031 31776 20076 31804
rect 20070 31764 20076 31776
rect 20128 31764 20134 31816
rect 20165 31807 20223 31813
rect 20165 31773 20177 31807
rect 20211 31804 20223 31807
rect 20346 31804 20352 31816
rect 20211 31776 20352 31804
rect 20211 31773 20223 31776
rect 20165 31767 20223 31773
rect 20346 31764 20352 31776
rect 20404 31764 20410 31816
rect 23198 31764 23204 31816
rect 23256 31804 23262 31816
rect 23293 31807 23351 31813
rect 23293 31804 23305 31807
rect 23256 31776 23305 31804
rect 23256 31764 23262 31776
rect 23293 31773 23305 31776
rect 23339 31773 23351 31807
rect 23293 31767 23351 31773
rect 23382 31764 23388 31816
rect 23440 31804 23446 31816
rect 24670 31804 24676 31816
rect 23440 31776 23485 31804
rect 24631 31776 24676 31804
rect 23440 31764 23446 31776
rect 24670 31764 24676 31776
rect 24728 31764 24734 31816
rect 26973 31807 27031 31813
rect 26973 31804 26985 31807
rect 26082 31776 26985 31804
rect 26973 31773 26985 31776
rect 27019 31773 27031 31807
rect 26973 31767 27031 31773
rect 27065 31807 27123 31813
rect 27065 31773 27077 31807
rect 27111 31804 27123 31807
rect 27614 31804 27620 31816
rect 27111 31776 27145 31804
rect 27575 31776 27620 31804
rect 27111 31773 27123 31776
rect 27065 31767 27123 31773
rect 15933 31739 15991 31745
rect 15933 31705 15945 31739
rect 15979 31736 15991 31739
rect 15979 31708 16013 31736
rect 15979 31705 15991 31708
rect 15933 31699 15991 31705
rect 1578 31668 1584 31680
rect 1539 31640 1584 31668
rect 1578 31628 1584 31640
rect 1636 31628 1642 31680
rect 6546 31628 6552 31680
rect 6604 31668 6610 31680
rect 6641 31671 6699 31677
rect 6641 31668 6653 31671
rect 6604 31640 6653 31668
rect 6604 31628 6610 31640
rect 6641 31637 6653 31640
rect 6687 31637 6699 31671
rect 8202 31668 8208 31680
rect 8163 31640 8208 31668
rect 6641 31631 6699 31637
rect 8202 31628 8208 31640
rect 8260 31628 8266 31680
rect 8294 31628 8300 31680
rect 8352 31668 8358 31680
rect 8352 31640 8397 31668
rect 8352 31628 8358 31640
rect 13998 31628 14004 31680
rect 14056 31668 14062 31680
rect 14645 31671 14703 31677
rect 14645 31668 14657 31671
rect 14056 31640 14657 31668
rect 14056 31628 14062 31640
rect 14645 31637 14657 31640
rect 14691 31637 14703 31671
rect 15562 31668 15568 31680
rect 15523 31640 15568 31668
rect 14645 31631 14703 31637
rect 15562 31628 15568 31640
rect 15620 31628 15626 31680
rect 16022 31668 16028 31680
rect 15983 31640 16028 31668
rect 16022 31628 16028 31640
rect 16080 31628 16086 31680
rect 17144 31668 17172 31764
rect 17402 31736 17408 31748
rect 17363 31708 17408 31736
rect 17402 31696 17408 31708
rect 17460 31696 17466 31748
rect 18708 31708 19564 31736
rect 17678 31668 17684 31680
rect 17144 31640 17684 31668
rect 17678 31628 17684 31640
rect 17736 31628 17742 31680
rect 17770 31628 17776 31680
rect 17828 31668 17834 31680
rect 18708 31668 18736 31708
rect 19426 31668 19432 31680
rect 17828 31640 18736 31668
rect 19387 31640 19432 31668
rect 17828 31628 17834 31640
rect 19426 31628 19432 31640
rect 19484 31628 19490 31680
rect 19536 31668 19564 31708
rect 21450 31696 21456 31748
rect 21508 31696 21514 31748
rect 26602 31696 26608 31748
rect 26660 31736 26666 31748
rect 27080 31736 27108 31767
rect 27614 31764 27620 31776
rect 27672 31764 27678 31816
rect 28074 31804 28080 31816
rect 28035 31776 28080 31804
rect 28074 31764 28080 31776
rect 28132 31764 28138 31816
rect 28537 31807 28595 31813
rect 28537 31773 28549 31807
rect 28583 31804 28595 31807
rect 28626 31804 28632 31816
rect 28583 31776 28632 31804
rect 28583 31773 28595 31776
rect 28537 31767 28595 31773
rect 28626 31764 28632 31776
rect 28684 31764 28690 31816
rect 28736 31813 28764 31912
rect 29086 31900 29092 31912
rect 29144 31900 29150 31952
rect 29362 31900 29368 31952
rect 29420 31940 29426 31952
rect 29420 31912 30052 31940
rect 29420 31900 29426 31912
rect 29181 31875 29239 31881
rect 29181 31841 29193 31875
rect 29227 31872 29239 31875
rect 29227 31844 29960 31872
rect 29227 31841 29239 31844
rect 29181 31835 29239 31841
rect 28721 31807 28779 31813
rect 28721 31773 28733 31807
rect 28767 31773 28779 31807
rect 28721 31767 28779 31773
rect 28813 31807 28871 31813
rect 28813 31773 28825 31807
rect 28859 31773 28871 31807
rect 28813 31767 28871 31773
rect 28905 31807 28963 31813
rect 28905 31773 28917 31807
rect 28951 31804 28963 31807
rect 28994 31804 29000 31816
rect 28951 31776 29000 31804
rect 28951 31773 28963 31776
rect 28905 31767 28963 31773
rect 26660 31708 27108 31736
rect 26660 31696 26666 31708
rect 28166 31696 28172 31748
rect 28224 31736 28230 31748
rect 28828 31736 28856 31767
rect 28994 31764 29000 31776
rect 29052 31764 29058 31816
rect 29546 31764 29552 31816
rect 29604 31804 29610 31816
rect 29932 31813 29960 31844
rect 30024 31813 30052 31912
rect 30742 31832 30748 31884
rect 30800 31872 30806 31884
rect 31297 31875 31355 31881
rect 31297 31872 31309 31875
rect 30800 31844 31309 31872
rect 30800 31832 30806 31844
rect 31297 31841 31309 31844
rect 31343 31872 31355 31875
rect 32766 31872 32772 31884
rect 31343 31844 32772 31872
rect 31343 31841 31355 31844
rect 31297 31835 31355 31841
rect 32766 31832 32772 31844
rect 32824 31832 32830 31884
rect 33318 31832 33324 31884
rect 33376 31872 33382 31884
rect 33376 31844 33824 31872
rect 33376 31832 33382 31844
rect 33796 31816 33824 31844
rect 29825 31807 29883 31813
rect 29825 31804 29837 31807
rect 29604 31776 29837 31804
rect 29604 31764 29610 31776
rect 29825 31773 29837 31776
rect 29871 31773 29883 31807
rect 29825 31767 29883 31773
rect 29917 31807 29975 31813
rect 29917 31773 29929 31807
rect 29963 31773 29975 31807
rect 29917 31767 29975 31773
rect 30009 31807 30067 31813
rect 30009 31773 30021 31807
rect 30055 31773 30067 31807
rect 30009 31767 30067 31773
rect 30193 31807 30251 31813
rect 30193 31773 30205 31807
rect 30239 31804 30251 31807
rect 30650 31804 30656 31816
rect 30239 31776 30656 31804
rect 30239 31773 30251 31776
rect 30193 31767 30251 31773
rect 30650 31764 30656 31776
rect 30708 31764 30714 31816
rect 30837 31807 30895 31813
rect 30837 31773 30849 31807
rect 30883 31804 30895 31807
rect 30926 31804 30932 31816
rect 30883 31776 30932 31804
rect 30883 31773 30895 31776
rect 30837 31767 30895 31773
rect 30926 31764 30932 31776
rect 30984 31764 30990 31816
rect 33689 31807 33747 31813
rect 33689 31804 33701 31807
rect 32706 31776 33701 31804
rect 33689 31773 33701 31776
rect 33735 31773 33747 31807
rect 33689 31767 33747 31773
rect 33778 31764 33784 31816
rect 33836 31804 33842 31816
rect 33836 31776 33881 31804
rect 33836 31764 33842 31776
rect 34514 31764 34520 31816
rect 34572 31804 34578 31816
rect 36909 31807 36967 31813
rect 36909 31804 36921 31807
rect 34572 31776 36921 31804
rect 34572 31764 34578 31776
rect 36909 31773 36921 31776
rect 36955 31773 36967 31807
rect 36909 31767 36967 31773
rect 31570 31736 31576 31748
rect 28224 31708 30880 31736
rect 31531 31708 31576 31736
rect 28224 31696 28230 31708
rect 26878 31668 26884 31680
rect 19536 31640 26884 31668
rect 26878 31628 26884 31640
rect 26936 31628 26942 31680
rect 27985 31671 28043 31677
rect 27985 31637 27997 31671
rect 28031 31668 28043 31671
rect 29730 31668 29736 31680
rect 28031 31640 29736 31668
rect 28031 31637 28043 31640
rect 27985 31631 28043 31637
rect 29730 31628 29736 31640
rect 29788 31628 29794 31680
rect 29914 31628 29920 31680
rect 29972 31668 29978 31680
rect 30745 31671 30803 31677
rect 30745 31668 30757 31671
rect 29972 31640 30757 31668
rect 29972 31628 29978 31640
rect 30745 31637 30757 31640
rect 30791 31637 30803 31671
rect 30852 31668 30880 31708
rect 31570 31696 31576 31708
rect 31628 31696 31634 31748
rect 32398 31668 32404 31680
rect 30852 31640 32404 31668
rect 30745 31631 30803 31637
rect 32398 31628 32404 31640
rect 32456 31628 32462 31680
rect 37090 31668 37096 31680
rect 37051 31640 37096 31668
rect 37090 31628 37096 31640
rect 37148 31628 37154 31680
rect 1104 31578 37628 31600
rect 1104 31526 4874 31578
rect 4926 31526 4938 31578
rect 4990 31526 5002 31578
rect 5054 31526 5066 31578
rect 5118 31526 5130 31578
rect 5182 31526 35594 31578
rect 35646 31526 35658 31578
rect 35710 31526 35722 31578
rect 35774 31526 35786 31578
rect 35838 31526 35850 31578
rect 35902 31526 37628 31578
rect 1104 31504 37628 31526
rect 7193 31467 7251 31473
rect 7193 31433 7205 31467
rect 7239 31433 7251 31467
rect 7193 31427 7251 31433
rect 7208 31396 7236 31427
rect 8938 31424 8944 31476
rect 8996 31464 9002 31476
rect 10413 31467 10471 31473
rect 10413 31464 10425 31467
rect 8996 31436 10425 31464
rect 8996 31424 9002 31436
rect 10413 31433 10425 31436
rect 10459 31433 10471 31467
rect 10413 31427 10471 31433
rect 10781 31467 10839 31473
rect 10781 31433 10793 31467
rect 10827 31464 10839 31467
rect 11698 31464 11704 31476
rect 10827 31436 11704 31464
rect 10827 31433 10839 31436
rect 10781 31427 10839 31433
rect 11698 31424 11704 31436
rect 11756 31424 11762 31476
rect 11885 31467 11943 31473
rect 11885 31433 11897 31467
rect 11931 31464 11943 31467
rect 17037 31467 17095 31473
rect 11931 31436 12434 31464
rect 11931 31433 11943 31436
rect 11885 31427 11943 31433
rect 7929 31399 7987 31405
rect 7929 31396 7941 31399
rect 7208 31368 7941 31396
rect 7929 31365 7941 31368
rect 7975 31365 7987 31399
rect 9214 31396 9220 31408
rect 9154 31368 9220 31396
rect 7929 31359 7987 31365
rect 9214 31356 9220 31368
rect 9272 31356 9278 31408
rect 10873 31399 10931 31405
rect 10873 31365 10885 31399
rect 10919 31396 10931 31399
rect 11514 31396 11520 31408
rect 10919 31368 11520 31396
rect 10919 31365 10931 31368
rect 10873 31359 10931 31365
rect 11514 31356 11520 31368
rect 11572 31356 11578 31408
rect 12406 31396 12434 31436
rect 17037 31433 17049 31467
rect 17083 31464 17095 31467
rect 17402 31464 17408 31476
rect 17083 31436 17408 31464
rect 17083 31433 17095 31436
rect 17037 31427 17095 31433
rect 17402 31424 17408 31436
rect 17460 31424 17466 31476
rect 17865 31467 17923 31473
rect 17865 31433 17877 31467
rect 17911 31464 17923 31467
rect 18693 31467 18751 31473
rect 18693 31464 18705 31467
rect 17911 31436 18705 31464
rect 17911 31433 17923 31436
rect 17865 31427 17923 31433
rect 18693 31433 18705 31436
rect 18739 31433 18751 31467
rect 19058 31464 19064 31476
rect 19019 31436 19064 31464
rect 18693 31427 18751 31433
rect 19058 31424 19064 31436
rect 19116 31424 19122 31476
rect 22833 31467 22891 31473
rect 22833 31433 22845 31467
rect 22879 31464 22891 31467
rect 23290 31464 23296 31476
rect 22879 31436 23296 31464
rect 22879 31433 22891 31436
rect 22833 31427 22891 31433
rect 23290 31424 23296 31436
rect 23348 31424 23354 31476
rect 24213 31467 24271 31473
rect 24213 31433 24225 31467
rect 24259 31433 24271 31467
rect 24213 31427 24271 31433
rect 14277 31399 14335 31405
rect 14277 31396 14289 31399
rect 12406 31368 14289 31396
rect 14277 31365 14289 31368
rect 14323 31365 14335 31399
rect 14277 31359 14335 31365
rect 15286 31356 15292 31408
rect 15344 31356 15350 31408
rect 16022 31356 16028 31408
rect 16080 31396 16086 31408
rect 17218 31396 17224 31408
rect 16080 31368 17224 31396
rect 16080 31356 16086 31368
rect 17218 31356 17224 31368
rect 17276 31396 17282 31408
rect 17770 31396 17776 31408
rect 17276 31368 17776 31396
rect 17276 31356 17282 31368
rect 17770 31356 17776 31368
rect 17828 31356 17834 31408
rect 24228 31396 24256 31427
rect 25038 31424 25044 31476
rect 25096 31464 25102 31476
rect 28994 31464 29000 31476
rect 25096 31436 29000 31464
rect 25096 31424 25102 31436
rect 24949 31399 25007 31405
rect 24949 31396 24961 31399
rect 17880 31368 22094 31396
rect 24228 31368 24961 31396
rect 17880 31340 17908 31368
rect 7006 31328 7012 31340
rect 6967 31300 7012 31328
rect 7006 31288 7012 31300
rect 7064 31288 7070 31340
rect 11701 31331 11759 31337
rect 11701 31297 11713 31331
rect 11747 31328 11759 31331
rect 11882 31328 11888 31340
rect 11747 31300 11888 31328
rect 11747 31297 11759 31300
rect 11701 31291 11759 31297
rect 11882 31288 11888 31300
rect 11940 31288 11946 31340
rect 11974 31288 11980 31340
rect 12032 31328 12038 31340
rect 12345 31331 12403 31337
rect 12345 31328 12357 31331
rect 12032 31300 12357 31328
rect 12032 31288 12038 31300
rect 12345 31297 12357 31300
rect 12391 31297 12403 31331
rect 12345 31291 12403 31297
rect 16853 31331 16911 31337
rect 16853 31297 16865 31331
rect 16899 31328 16911 31331
rect 16899 31300 17540 31328
rect 16899 31297 16911 31300
rect 16853 31291 16911 31297
rect 6454 31220 6460 31272
rect 6512 31260 6518 31272
rect 7653 31263 7711 31269
rect 7653 31260 7665 31263
rect 6512 31232 7665 31260
rect 6512 31220 6518 31232
rect 7653 31229 7665 31232
rect 7699 31229 7711 31263
rect 7653 31223 7711 31229
rect 10870 31220 10876 31272
rect 10928 31260 10934 31272
rect 10965 31263 11023 31269
rect 10965 31260 10977 31263
rect 10928 31232 10977 31260
rect 10928 31220 10934 31232
rect 10965 31229 10977 31232
rect 11011 31229 11023 31263
rect 10965 31223 11023 31229
rect 12250 31220 12256 31272
rect 12308 31260 12314 31272
rect 13173 31263 13231 31269
rect 13173 31260 13185 31263
rect 12308 31232 13185 31260
rect 12308 31220 12314 31232
rect 13173 31229 13185 31232
rect 13219 31260 13231 31263
rect 13814 31260 13820 31272
rect 13219 31232 13820 31260
rect 13219 31229 13231 31232
rect 13173 31223 13231 31229
rect 13814 31220 13820 31232
rect 13872 31260 13878 31272
rect 14001 31263 14059 31269
rect 14001 31260 14013 31263
rect 13872 31232 14013 31260
rect 13872 31220 13878 31232
rect 14001 31229 14013 31232
rect 14047 31229 14059 31263
rect 14001 31223 14059 31229
rect 17512 31201 17540 31300
rect 17862 31288 17868 31340
rect 17920 31288 17926 31340
rect 17957 31331 18015 31337
rect 17957 31297 17969 31331
rect 18003 31328 18015 31331
rect 19886 31328 19892 31340
rect 18003 31300 19892 31328
rect 18003 31297 18015 31300
rect 17957 31291 18015 31297
rect 19886 31288 19892 31300
rect 19944 31288 19950 31340
rect 20717 31331 20775 31337
rect 20717 31297 20729 31331
rect 20763 31328 20775 31331
rect 20898 31328 20904 31340
rect 20763 31300 20904 31328
rect 20763 31297 20775 31300
rect 20717 31291 20775 31297
rect 20898 31288 20904 31300
rect 20956 31288 20962 31340
rect 21266 31328 21272 31340
rect 21227 31300 21272 31328
rect 21266 31288 21272 31300
rect 21324 31288 21330 31340
rect 18141 31263 18199 31269
rect 18141 31229 18153 31263
rect 18187 31229 18199 31263
rect 19150 31260 19156 31272
rect 19111 31232 19156 31260
rect 18141 31223 18199 31229
rect 17497 31195 17555 31201
rect 17497 31161 17509 31195
rect 17543 31161 17555 31195
rect 17497 31155 17555 31161
rect 18156 31192 18184 31223
rect 19150 31220 19156 31232
rect 19208 31220 19214 31272
rect 19334 31260 19340 31272
rect 19295 31232 19340 31260
rect 19334 31220 19340 31232
rect 19392 31220 19398 31272
rect 20441 31195 20499 31201
rect 20441 31192 20453 31195
rect 18156 31164 20453 31192
rect 9398 31124 9404 31136
rect 9359 31096 9404 31124
rect 9398 31084 9404 31096
rect 9456 31084 9462 31136
rect 15749 31127 15807 31133
rect 15749 31093 15761 31127
rect 15795 31124 15807 31127
rect 16574 31124 16580 31136
rect 15795 31096 16580 31124
rect 15795 31093 15807 31096
rect 15749 31087 15807 31093
rect 16574 31084 16580 31096
rect 16632 31084 16638 31136
rect 17954 31084 17960 31136
rect 18012 31124 18018 31136
rect 18156 31124 18184 31164
rect 20441 31161 20453 31164
rect 20487 31161 20499 31195
rect 22066 31192 22094 31368
rect 24949 31365 24961 31368
rect 24995 31365 25007 31399
rect 26418 31396 26424 31408
rect 26174 31368 26424 31396
rect 24949 31359 25007 31365
rect 26418 31356 26424 31368
rect 26476 31356 26482 31408
rect 22741 31331 22799 31337
rect 22741 31297 22753 31331
rect 22787 31328 22799 31331
rect 23842 31328 23848 31340
rect 22787 31300 23848 31328
rect 22787 31297 22799 31300
rect 22741 31291 22799 31297
rect 23842 31288 23848 31300
rect 23900 31288 23906 31340
rect 24029 31331 24087 31337
rect 24029 31297 24041 31331
rect 24075 31328 24087 31331
rect 24578 31328 24584 31340
rect 24075 31300 24584 31328
rect 24075 31297 24087 31300
rect 24029 31291 24087 31297
rect 24578 31288 24584 31300
rect 24636 31288 24642 31340
rect 22646 31260 22652 31272
rect 22607 31232 22652 31260
rect 22646 31220 22652 31232
rect 22704 31220 22710 31272
rect 22922 31220 22928 31272
rect 22980 31260 22986 31272
rect 24670 31260 24676 31272
rect 22980 31232 24676 31260
rect 22980 31220 22986 31232
rect 24670 31220 24676 31232
rect 24728 31220 24734 31272
rect 26421 31195 26479 31201
rect 22066 31164 23704 31192
rect 20441 31155 20499 31161
rect 21358 31124 21364 31136
rect 18012 31096 18184 31124
rect 21319 31096 21364 31124
rect 18012 31084 18018 31096
rect 21358 31084 21364 31096
rect 21416 31084 21422 31136
rect 23201 31127 23259 31133
rect 23201 31093 23213 31127
rect 23247 31124 23259 31127
rect 23566 31124 23572 31136
rect 23247 31096 23572 31124
rect 23247 31093 23259 31096
rect 23201 31087 23259 31093
rect 23566 31084 23572 31096
rect 23624 31084 23630 31136
rect 23676 31124 23704 31164
rect 26421 31161 26433 31195
rect 26467 31192 26479 31195
rect 26804 31192 26832 31436
rect 28994 31424 29000 31436
rect 29052 31424 29058 31476
rect 33594 31464 33600 31476
rect 30392 31436 33600 31464
rect 26878 31356 26884 31408
rect 26936 31396 26942 31408
rect 30392 31405 30420 31436
rect 33594 31424 33600 31436
rect 33652 31424 33658 31476
rect 33781 31467 33839 31473
rect 33781 31433 33793 31467
rect 33827 31464 33839 31467
rect 34514 31464 34520 31476
rect 33827 31436 34520 31464
rect 33827 31433 33839 31436
rect 33781 31427 33839 31433
rect 34514 31424 34520 31436
rect 34572 31424 34578 31476
rect 34609 31467 34667 31473
rect 34609 31433 34621 31467
rect 34655 31464 34667 31467
rect 36906 31464 36912 31476
rect 34655 31436 36912 31464
rect 34655 31433 34667 31436
rect 34609 31427 34667 31433
rect 36906 31424 36912 31436
rect 36964 31424 36970 31476
rect 30377 31399 30435 31405
rect 26936 31368 28120 31396
rect 26936 31356 26942 31368
rect 27982 31328 27988 31340
rect 27943 31300 27988 31328
rect 27982 31288 27988 31300
rect 28040 31288 28046 31340
rect 28092 31328 28120 31368
rect 30377 31365 30389 31399
rect 30423 31365 30435 31399
rect 30377 31359 30435 31365
rect 31005 31399 31063 31405
rect 31005 31365 31017 31399
rect 31051 31396 31063 31399
rect 31110 31396 31116 31408
rect 31051 31368 31116 31396
rect 31051 31365 31063 31368
rect 31005 31359 31063 31365
rect 31110 31356 31116 31368
rect 31168 31356 31174 31408
rect 31205 31399 31263 31405
rect 31205 31365 31217 31399
rect 31251 31396 31263 31399
rect 31294 31396 31300 31408
rect 31251 31368 31300 31396
rect 31251 31365 31263 31368
rect 31205 31359 31263 31365
rect 31294 31356 31300 31368
rect 31352 31396 31358 31408
rect 31478 31396 31484 31408
rect 31352 31368 31484 31396
rect 31352 31356 31358 31368
rect 31478 31356 31484 31368
rect 31536 31356 31542 31408
rect 31662 31356 31668 31408
rect 31720 31396 31726 31408
rect 32677 31399 32735 31405
rect 32677 31396 32689 31399
rect 31720 31368 32689 31396
rect 31720 31356 31726 31368
rect 32677 31365 32689 31368
rect 32723 31365 32735 31399
rect 32677 31359 32735 31365
rect 32585 31331 32643 31337
rect 32585 31328 32597 31331
rect 28092 31300 32597 31328
rect 32585 31297 32597 31300
rect 32631 31297 32643 31331
rect 33597 31331 33655 31337
rect 33597 31328 33609 31331
rect 32585 31291 32643 31297
rect 33060 31300 33609 31328
rect 32401 31263 32459 31269
rect 32401 31260 32413 31263
rect 26467 31164 26832 31192
rect 26896 31232 32413 31260
rect 26467 31161 26479 31164
rect 26421 31155 26479 31161
rect 26896 31124 26924 31232
rect 32401 31229 32413 31232
rect 32447 31229 32459 31263
rect 32401 31223 32459 31229
rect 27525 31195 27583 31201
rect 27525 31161 27537 31195
rect 27571 31192 27583 31195
rect 27614 31192 27620 31204
rect 27571 31164 27620 31192
rect 27571 31161 27583 31164
rect 27525 31155 27583 31161
rect 27614 31152 27620 31164
rect 27672 31192 27678 31204
rect 29270 31192 29276 31204
rect 27672 31164 29276 31192
rect 27672 31152 27678 31164
rect 29270 31152 29276 31164
rect 29328 31152 29334 31204
rect 30834 31192 30840 31204
rect 30795 31164 30840 31192
rect 30834 31152 30840 31164
rect 30892 31152 30898 31204
rect 27890 31124 27896 31136
rect 23676 31096 26924 31124
rect 27803 31096 27896 31124
rect 27890 31084 27896 31096
rect 27948 31124 27954 31136
rect 28442 31124 28448 31136
rect 27948 31096 28448 31124
rect 27948 31084 27954 31096
rect 28442 31084 28448 31096
rect 28500 31084 28506 31136
rect 29089 31127 29147 31133
rect 29089 31093 29101 31127
rect 29135 31124 29147 31127
rect 30742 31124 30748 31136
rect 29135 31096 30748 31124
rect 29135 31093 29147 31096
rect 29089 31087 29147 31093
rect 30742 31084 30748 31096
rect 30800 31084 30806 31136
rect 30926 31084 30932 31136
rect 30984 31124 30990 31136
rect 31021 31127 31079 31133
rect 31021 31124 31033 31127
rect 30984 31096 31033 31124
rect 30984 31084 30990 31096
rect 31021 31093 31033 31096
rect 31067 31093 31079 31127
rect 32416 31124 32444 31223
rect 33060 31201 33088 31300
rect 33597 31297 33609 31300
rect 33643 31297 33655 31331
rect 33597 31291 33655 31297
rect 34330 31288 34336 31340
rect 34388 31328 34394 31340
rect 34425 31331 34483 31337
rect 34425 31328 34437 31331
rect 34388 31300 34437 31328
rect 34388 31288 34394 31300
rect 34425 31297 34437 31300
rect 34471 31297 34483 31331
rect 34425 31291 34483 31297
rect 33045 31195 33103 31201
rect 33045 31161 33057 31195
rect 33091 31161 33103 31195
rect 33045 31155 33103 31161
rect 33594 31124 33600 31136
rect 32416 31096 33600 31124
rect 31021 31087 31079 31093
rect 33594 31084 33600 31096
rect 33652 31084 33658 31136
rect 1104 31034 37628 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 37628 31034
rect 1104 30960 37628 30982
rect 8202 30920 8208 30932
rect 8163 30892 8208 30920
rect 8202 30880 8208 30892
rect 8260 30880 8266 30932
rect 10962 30880 10968 30932
rect 11020 30920 11026 30932
rect 11793 30923 11851 30929
rect 11793 30920 11805 30923
rect 11020 30892 11805 30920
rect 11020 30880 11026 30892
rect 11793 30889 11805 30892
rect 11839 30889 11851 30923
rect 11793 30883 11851 30889
rect 11882 30880 11888 30932
rect 11940 30920 11946 30932
rect 14737 30923 14795 30929
rect 14737 30920 14749 30923
rect 11940 30892 14749 30920
rect 11940 30880 11946 30892
rect 14737 30889 14749 30892
rect 14783 30889 14795 30923
rect 14737 30883 14795 30889
rect 15933 30923 15991 30929
rect 15933 30889 15945 30923
rect 15979 30920 15991 30923
rect 16022 30920 16028 30932
rect 15979 30892 16028 30920
rect 15979 30889 15991 30892
rect 15933 30883 15991 30889
rect 16022 30880 16028 30892
rect 16080 30880 16086 30932
rect 16114 30880 16120 30932
rect 16172 30920 16178 30932
rect 19334 30920 19340 30932
rect 16172 30892 19340 30920
rect 16172 30880 16178 30892
rect 19334 30880 19340 30892
rect 19392 30880 19398 30932
rect 19429 30923 19487 30929
rect 19429 30889 19441 30923
rect 19475 30920 19487 30923
rect 19610 30920 19616 30932
rect 19475 30892 19616 30920
rect 19475 30889 19487 30892
rect 19429 30883 19487 30889
rect 19610 30880 19616 30892
rect 19668 30880 19674 30932
rect 21177 30923 21235 30929
rect 21177 30889 21189 30923
rect 21223 30920 21235 30923
rect 23842 30920 23848 30932
rect 21223 30892 23848 30920
rect 21223 30889 21235 30892
rect 21177 30883 21235 30889
rect 23842 30880 23848 30892
rect 23900 30880 23906 30932
rect 24578 30920 24584 30932
rect 24539 30892 24584 30920
rect 24578 30880 24584 30892
rect 24636 30880 24642 30932
rect 27982 30880 27988 30932
rect 28040 30920 28046 30932
rect 28721 30923 28779 30929
rect 28721 30920 28733 30923
rect 28040 30892 28733 30920
rect 28040 30880 28046 30892
rect 28721 30889 28733 30892
rect 28767 30920 28779 30923
rect 29730 30920 29736 30932
rect 28767 30892 29592 30920
rect 29691 30892 29736 30920
rect 28767 30889 28779 30892
rect 28721 30883 28779 30889
rect 12618 30812 12624 30864
rect 12676 30852 12682 30864
rect 13357 30855 13415 30861
rect 13357 30852 13369 30855
rect 12676 30824 13369 30852
rect 12676 30812 12682 30824
rect 13357 30821 13369 30824
rect 13403 30821 13415 30855
rect 13357 30815 13415 30821
rect 15102 30812 15108 30864
rect 15160 30812 15166 30864
rect 21266 30852 21272 30864
rect 18708 30824 21272 30852
rect 7098 30784 7104 30796
rect 6472 30756 7104 30784
rect 6472 30728 6500 30756
rect 7098 30744 7104 30756
rect 7156 30744 7162 30796
rect 9766 30744 9772 30796
rect 9824 30784 9830 30796
rect 9953 30787 10011 30793
rect 9953 30784 9965 30787
rect 9824 30756 9965 30784
rect 9824 30744 9830 30756
rect 9953 30753 9965 30756
rect 9999 30753 10011 30787
rect 9953 30747 10011 30753
rect 11514 30744 11520 30796
rect 11572 30784 11578 30796
rect 12253 30787 12311 30793
rect 12253 30784 12265 30787
rect 11572 30756 12265 30784
rect 11572 30744 11578 30756
rect 12253 30753 12265 30756
rect 12299 30753 12311 30787
rect 12253 30747 12311 30753
rect 12345 30787 12403 30793
rect 12345 30753 12357 30787
rect 12391 30784 12403 30787
rect 12526 30784 12532 30796
rect 12391 30756 12532 30784
rect 12391 30753 12403 30756
rect 12345 30747 12403 30753
rect 12526 30744 12532 30756
rect 12584 30744 12590 30796
rect 14826 30744 14832 30796
rect 14884 30784 14890 30796
rect 15120 30784 15148 30812
rect 15289 30787 15347 30793
rect 15289 30784 15301 30787
rect 14884 30756 15301 30784
rect 14884 30744 14890 30756
rect 15289 30753 15301 30756
rect 15335 30753 15347 30787
rect 15289 30747 15347 30753
rect 17310 30744 17316 30796
rect 17368 30784 17374 30796
rect 18708 30793 18736 30824
rect 21266 30812 21272 30824
rect 21324 30812 21330 30864
rect 28074 30812 28080 30864
rect 28132 30852 28138 30864
rect 28902 30852 28908 30864
rect 28132 30824 28908 30852
rect 28132 30812 28138 30824
rect 28902 30812 28908 30824
rect 28960 30812 28966 30864
rect 29564 30852 29592 30892
rect 29730 30880 29736 30892
rect 29788 30880 29794 30932
rect 30101 30923 30159 30929
rect 30101 30889 30113 30923
rect 30147 30920 30159 30923
rect 30558 30920 30564 30932
rect 30147 30892 30564 30920
rect 30147 30889 30159 30892
rect 30101 30883 30159 30889
rect 30558 30880 30564 30892
rect 30616 30920 30622 30932
rect 31202 30920 31208 30932
rect 30616 30892 31208 30920
rect 30616 30880 30622 30892
rect 31202 30880 31208 30892
rect 31260 30920 31266 30932
rect 32677 30923 32735 30929
rect 32677 30920 32689 30923
rect 31260 30892 32689 30920
rect 31260 30880 31266 30892
rect 32677 30889 32689 30892
rect 32723 30889 32735 30923
rect 34330 30920 34336 30932
rect 34291 30892 34336 30920
rect 32677 30883 32735 30889
rect 34330 30880 34336 30892
rect 34388 30880 34394 30932
rect 30834 30852 30840 30864
rect 29564 30824 30840 30852
rect 30834 30812 30840 30824
rect 30892 30812 30898 30864
rect 17405 30787 17463 30793
rect 17405 30784 17417 30787
rect 17368 30756 17417 30784
rect 17368 30744 17374 30756
rect 17405 30753 17417 30756
rect 17451 30753 17463 30787
rect 17405 30747 17463 30753
rect 18693 30787 18751 30793
rect 18693 30753 18705 30787
rect 18739 30753 18751 30787
rect 19886 30784 19892 30796
rect 19847 30756 19892 30784
rect 18693 30747 18751 30753
rect 19886 30744 19892 30756
rect 19944 30744 19950 30796
rect 19978 30744 19984 30796
rect 20036 30784 20042 30796
rect 20036 30756 20081 30784
rect 20036 30744 20042 30756
rect 22186 30744 22192 30796
rect 22244 30784 22250 30796
rect 22244 30756 22968 30784
rect 22244 30744 22250 30756
rect 22940 30728 22968 30756
rect 24854 30744 24860 30796
rect 24912 30784 24918 30796
rect 25130 30784 25136 30796
rect 24912 30756 25136 30784
rect 24912 30744 24918 30756
rect 25130 30744 25136 30756
rect 25188 30744 25194 30796
rect 29914 30784 29920 30796
rect 27632 30756 29920 30784
rect 27632 30728 27660 30756
rect 29914 30744 29920 30756
rect 29972 30744 29978 30796
rect 30742 30744 30748 30796
rect 30800 30784 30806 30796
rect 30929 30787 30987 30793
rect 30929 30784 30941 30787
rect 30800 30756 30941 30784
rect 30800 30744 30806 30756
rect 30929 30753 30941 30756
rect 30975 30753 30987 30787
rect 30929 30747 30987 30753
rect 31205 30787 31263 30793
rect 31205 30753 31217 30787
rect 31251 30784 31263 30787
rect 32398 30784 32404 30796
rect 31251 30756 32404 30784
rect 31251 30753 31263 30756
rect 31205 30747 31263 30753
rect 32398 30744 32404 30756
rect 32456 30744 32462 30796
rect 33594 30744 33600 30796
rect 33652 30784 33658 30796
rect 33689 30787 33747 30793
rect 33689 30784 33701 30787
rect 33652 30756 33701 30784
rect 33652 30744 33658 30756
rect 33689 30753 33701 30756
rect 33735 30753 33747 30787
rect 33689 30747 33747 30753
rect 6454 30716 6460 30728
rect 6415 30688 6460 30716
rect 6454 30676 6460 30688
rect 6512 30676 6518 30728
rect 9214 30716 9220 30728
rect 9175 30688 9220 30716
rect 9214 30676 9220 30688
rect 9272 30676 9278 30728
rect 12158 30716 12164 30728
rect 12119 30688 12164 30716
rect 12158 30676 12164 30688
rect 12216 30676 12222 30728
rect 15105 30719 15163 30725
rect 15105 30685 15117 30719
rect 15151 30716 15163 30719
rect 15562 30716 15568 30728
rect 15151 30688 15568 30716
rect 15151 30685 15163 30688
rect 15105 30679 15163 30685
rect 15562 30676 15568 30688
rect 15620 30676 15626 30728
rect 17678 30676 17684 30728
rect 17736 30716 17742 30728
rect 17736 30688 17781 30716
rect 17736 30676 17742 30688
rect 18506 30676 18512 30728
rect 18564 30716 18570 30728
rect 18877 30719 18935 30725
rect 18877 30716 18889 30719
rect 18564 30688 18889 30716
rect 18564 30676 18570 30688
rect 18877 30685 18889 30688
rect 18923 30685 18935 30719
rect 18877 30679 18935 30685
rect 19150 30676 19156 30728
rect 19208 30716 19214 30728
rect 19797 30719 19855 30725
rect 19797 30716 19809 30719
rect 19208 30688 19809 30716
rect 19208 30676 19214 30688
rect 19797 30685 19809 30688
rect 19843 30716 19855 30719
rect 20806 30716 20812 30728
rect 19843 30688 20812 30716
rect 19843 30685 19855 30688
rect 19797 30679 19855 30685
rect 20806 30676 20812 30688
rect 20864 30676 20870 30728
rect 22922 30676 22928 30728
rect 22980 30716 22986 30728
rect 23566 30716 23572 30728
rect 22980 30688 23025 30716
rect 23527 30688 23572 30716
rect 22980 30676 22986 30688
rect 23566 30676 23572 30688
rect 23624 30676 23630 30728
rect 24946 30716 24952 30728
rect 24907 30688 24952 30716
rect 24946 30676 24952 30688
rect 25004 30676 25010 30728
rect 25958 30716 25964 30728
rect 25919 30688 25964 30716
rect 25958 30676 25964 30688
rect 26016 30676 26022 30728
rect 26602 30716 26608 30728
rect 26563 30688 26608 30716
rect 26602 30676 26608 30688
rect 26660 30676 26666 30728
rect 27338 30716 27344 30728
rect 27299 30688 27344 30716
rect 27338 30676 27344 30688
rect 27396 30676 27402 30728
rect 27434 30719 27492 30725
rect 27434 30685 27446 30719
rect 27480 30685 27492 30719
rect 27434 30679 27492 30685
rect 6638 30608 6644 30660
rect 6696 30648 6702 30660
rect 6733 30651 6791 30657
rect 6733 30648 6745 30651
rect 6696 30620 6745 30648
rect 6696 30608 6702 30620
rect 6733 30617 6745 30620
rect 6779 30617 6791 30651
rect 10781 30651 10839 30657
rect 6733 30611 6791 30617
rect 6886 30620 7222 30648
rect 6546 30540 6552 30592
rect 6604 30580 6610 30592
rect 6886 30580 6914 30620
rect 10781 30617 10793 30651
rect 10827 30648 10839 30651
rect 11974 30648 11980 30660
rect 10827 30620 11980 30648
rect 10827 30617 10839 30620
rect 10781 30611 10839 30617
rect 11974 30608 11980 30620
rect 12032 30608 12038 30660
rect 13630 30648 13636 30660
rect 13591 30620 13636 30648
rect 13630 30608 13636 30620
rect 13688 30608 13694 30660
rect 15197 30651 15255 30657
rect 15197 30617 15209 30651
rect 15243 30648 15255 30651
rect 15243 30620 16160 30648
rect 15243 30617 15255 30620
rect 15197 30611 15255 30617
rect 9306 30580 9312 30592
rect 6604 30552 6914 30580
rect 9267 30552 9312 30580
rect 6604 30540 6610 30552
rect 9306 30540 9312 30552
rect 9364 30540 9370 30592
rect 16132 30580 16160 30620
rect 16390 30608 16396 30660
rect 16448 30608 16454 30660
rect 21358 30608 21364 30660
rect 21416 30648 21422 30660
rect 22649 30651 22707 30657
rect 21416 30620 21482 30648
rect 21416 30608 21422 30620
rect 22649 30617 22661 30651
rect 22695 30648 22707 30651
rect 22695 30620 23428 30648
rect 22695 30617 22707 30620
rect 22649 30611 22707 30617
rect 16574 30580 16580 30592
rect 16132 30552 16580 30580
rect 16574 30540 16580 30552
rect 16632 30540 16638 30592
rect 23400 30589 23428 30620
rect 23842 30608 23848 30660
rect 23900 30648 23906 30660
rect 25041 30651 25099 30657
rect 25041 30648 25053 30651
rect 23900 30620 25053 30648
rect 23900 30608 23906 30620
rect 25041 30617 25053 30620
rect 25087 30617 25099 30651
rect 25041 30611 25099 30617
rect 27246 30608 27252 30660
rect 27304 30648 27310 30660
rect 27448 30648 27476 30679
rect 27614 30676 27620 30728
rect 27672 30716 27678 30728
rect 27890 30725 27896 30728
rect 27847 30719 27896 30725
rect 27672 30688 27765 30716
rect 27672 30676 27678 30688
rect 27847 30685 27859 30719
rect 27893 30685 27896 30719
rect 27847 30679 27896 30685
rect 27890 30676 27896 30679
rect 27948 30676 27954 30728
rect 27982 30676 27988 30728
rect 28040 30676 28046 30728
rect 28442 30716 28448 30728
rect 28403 30688 28448 30716
rect 28442 30676 28448 30688
rect 28500 30676 28506 30728
rect 28994 30676 29000 30728
rect 29052 30716 29058 30728
rect 30193 30719 30251 30725
rect 30193 30716 30205 30719
rect 29052 30688 30205 30716
rect 29052 30676 29058 30688
rect 30193 30685 30205 30688
rect 30239 30685 30251 30719
rect 30193 30679 30251 30685
rect 27304 30620 27476 30648
rect 27709 30651 27767 30657
rect 27304 30608 27310 30620
rect 27709 30617 27721 30651
rect 27755 30648 27767 30651
rect 28000 30648 28028 30676
rect 33686 30648 33692 30660
rect 27755 30620 28028 30648
rect 32430 30620 33692 30648
rect 27755 30617 27767 30620
rect 27709 30611 27767 30617
rect 33686 30608 33692 30620
rect 33744 30608 33750 30660
rect 23385 30583 23443 30589
rect 23385 30549 23397 30583
rect 23431 30549 23443 30583
rect 23385 30543 23443 30549
rect 25222 30540 25228 30592
rect 25280 30580 25286 30592
rect 25777 30583 25835 30589
rect 25777 30580 25789 30583
rect 25280 30552 25789 30580
rect 25280 30540 25286 30552
rect 25777 30549 25789 30552
rect 25823 30549 25835 30583
rect 26510 30580 26516 30592
rect 26471 30552 26516 30580
rect 25777 30543 25835 30549
rect 26510 30540 26516 30552
rect 26568 30540 26574 30592
rect 27798 30540 27804 30592
rect 27856 30580 27862 30592
rect 27985 30583 28043 30589
rect 27985 30580 27997 30583
rect 27856 30552 27997 30580
rect 27856 30540 27862 30552
rect 27985 30549 27997 30552
rect 28031 30549 28043 30583
rect 27985 30543 28043 30549
rect 28442 30540 28448 30592
rect 28500 30580 28506 30592
rect 33873 30583 33931 30589
rect 33873 30580 33885 30583
rect 28500 30552 33885 30580
rect 28500 30540 28506 30552
rect 33873 30549 33885 30552
rect 33919 30549 33931 30583
rect 33873 30543 33931 30549
rect 33962 30540 33968 30592
rect 34020 30580 34026 30592
rect 34020 30552 34065 30580
rect 34020 30540 34026 30552
rect 1104 30490 37628 30512
rect 1104 30438 4874 30490
rect 4926 30438 4938 30490
rect 4990 30438 5002 30490
rect 5054 30438 5066 30490
rect 5118 30438 5130 30490
rect 5182 30438 35594 30490
rect 35646 30438 35658 30490
rect 35710 30438 35722 30490
rect 35774 30438 35786 30490
rect 35838 30438 35850 30490
rect 35902 30438 37628 30490
rect 1104 30416 37628 30438
rect 8294 30376 8300 30388
rect 8128 30348 8300 30376
rect 7285 30311 7343 30317
rect 7285 30277 7297 30311
rect 7331 30308 7343 30311
rect 8128 30308 8156 30348
rect 8294 30336 8300 30348
rect 8352 30376 8358 30388
rect 9398 30376 9404 30388
rect 8352 30348 9404 30376
rect 8352 30336 8358 30348
rect 9398 30336 9404 30348
rect 9456 30376 9462 30388
rect 9585 30379 9643 30385
rect 9585 30376 9597 30379
rect 9456 30348 9597 30376
rect 9456 30336 9462 30348
rect 9585 30345 9597 30348
rect 9631 30345 9643 30379
rect 9585 30339 9643 30345
rect 11146 30336 11152 30388
rect 11204 30376 11210 30388
rect 12526 30376 12532 30388
rect 11204 30348 12532 30376
rect 11204 30336 11210 30348
rect 12526 30336 12532 30348
rect 12584 30336 12590 30388
rect 16574 30336 16580 30388
rect 16632 30376 16638 30388
rect 19058 30376 19064 30388
rect 16632 30348 19064 30376
rect 16632 30336 16638 30348
rect 7331 30280 8156 30308
rect 7331 30277 7343 30280
rect 7285 30271 7343 30277
rect 8202 30268 8208 30320
rect 8260 30308 8266 30320
rect 8481 30311 8539 30317
rect 8481 30308 8493 30311
rect 8260 30280 8493 30308
rect 8260 30268 8266 30280
rect 8481 30277 8493 30280
rect 8527 30277 8539 30311
rect 8481 30271 8539 30277
rect 9493 30311 9551 30317
rect 9493 30277 9505 30311
rect 9539 30308 9551 30311
rect 10781 30311 10839 30317
rect 10781 30308 10793 30311
rect 9539 30280 10793 30308
rect 9539 30277 9551 30280
rect 9493 30271 9551 30277
rect 10781 30277 10793 30280
rect 10827 30308 10839 30311
rect 12894 30308 12900 30320
rect 10827 30280 12900 30308
rect 10827 30277 10839 30280
rect 10781 30271 10839 30277
rect 12894 30268 12900 30280
rect 12952 30308 12958 30320
rect 13265 30311 13323 30317
rect 13265 30308 13277 30311
rect 12952 30280 13277 30308
rect 12952 30268 12958 30280
rect 13265 30277 13277 30280
rect 13311 30277 13323 30311
rect 14826 30308 14832 30320
rect 14787 30280 14832 30308
rect 13265 30271 13323 30277
rect 14826 30268 14832 30280
rect 14884 30268 14890 30320
rect 16209 30311 16267 30317
rect 16209 30277 16221 30311
rect 16255 30308 16267 30311
rect 16390 30308 16396 30320
rect 16255 30280 16396 30308
rect 16255 30277 16267 30280
rect 16209 30271 16267 30277
rect 16390 30268 16396 30280
rect 16448 30268 16454 30320
rect 17218 30308 17224 30320
rect 17179 30280 17224 30308
rect 17218 30268 17224 30280
rect 17276 30268 17282 30320
rect 17328 30317 17356 30348
rect 19058 30336 19064 30348
rect 19116 30336 19122 30388
rect 25409 30379 25467 30385
rect 22112 30348 22416 30376
rect 17313 30311 17371 30317
rect 17313 30277 17325 30311
rect 17359 30277 17371 30311
rect 17313 30271 17371 30277
rect 17678 30268 17684 30320
rect 17736 30308 17742 30320
rect 19337 30311 19395 30317
rect 17736 30280 19104 30308
rect 17736 30268 17742 30280
rect 7193 30243 7251 30249
rect 7193 30209 7205 30243
rect 7239 30209 7251 30243
rect 7193 30203 7251 30209
rect 6825 30107 6883 30113
rect 6825 30073 6837 30107
rect 6871 30104 6883 30107
rect 7006 30104 7012 30116
rect 6871 30076 7012 30104
rect 6871 30073 6883 30076
rect 6825 30067 6883 30073
rect 7006 30064 7012 30076
rect 7064 30064 7070 30116
rect 7208 30104 7236 30203
rect 8294 30200 8300 30252
rect 8352 30240 8358 30252
rect 8389 30243 8447 30249
rect 8389 30240 8401 30243
rect 8352 30212 8401 30240
rect 8352 30200 8358 30212
rect 8389 30209 8401 30212
rect 8435 30209 8447 30243
rect 8389 30203 8447 30209
rect 10873 30243 10931 30249
rect 10873 30209 10885 30243
rect 10919 30240 10931 30243
rect 11238 30240 11244 30252
rect 10919 30212 11244 30240
rect 10919 30209 10931 30212
rect 10873 30203 10931 30209
rect 11238 30200 11244 30212
rect 11296 30240 11302 30252
rect 12066 30240 12072 30252
rect 11296 30212 12072 30240
rect 11296 30200 11302 30212
rect 12066 30200 12072 30212
rect 12124 30200 12130 30252
rect 12345 30243 12403 30249
rect 12345 30209 12357 30243
rect 12391 30209 12403 30243
rect 12345 30203 12403 30209
rect 7469 30175 7527 30181
rect 7469 30141 7481 30175
rect 7515 30172 7527 30175
rect 8202 30172 8208 30184
rect 7515 30144 8208 30172
rect 7515 30141 7527 30144
rect 7469 30135 7527 30141
rect 8202 30132 8208 30144
rect 8260 30132 8266 30184
rect 8665 30175 8723 30181
rect 8665 30141 8677 30175
rect 8711 30172 8723 30175
rect 9401 30175 9459 30181
rect 9401 30172 9413 30175
rect 8711 30144 9413 30172
rect 8711 30141 8723 30144
rect 8665 30135 8723 30141
rect 9401 30141 9413 30144
rect 9447 30172 9459 30175
rect 9582 30172 9588 30184
rect 9447 30144 9588 30172
rect 9447 30141 9459 30144
rect 9401 30135 9459 30141
rect 9582 30132 9588 30144
rect 9640 30132 9646 30184
rect 10965 30175 11023 30181
rect 10965 30141 10977 30175
rect 11011 30172 11023 30175
rect 11146 30172 11152 30184
rect 11011 30144 11152 30172
rect 11011 30141 11023 30144
rect 10965 30135 11023 30141
rect 11146 30132 11152 30144
rect 11204 30132 11210 30184
rect 12161 30175 12219 30181
rect 12161 30141 12173 30175
rect 12207 30172 12219 30175
rect 12250 30172 12256 30184
rect 12207 30144 12256 30172
rect 12207 30141 12219 30144
rect 12161 30135 12219 30141
rect 12250 30132 12256 30144
rect 12308 30132 12314 30184
rect 8021 30107 8079 30113
rect 8021 30104 8033 30107
rect 7208 30076 8033 30104
rect 8021 30073 8033 30076
rect 8067 30073 8079 30107
rect 8021 30067 8079 30073
rect 9122 30064 9128 30116
rect 9180 30104 9186 30116
rect 10413 30107 10471 30113
rect 10413 30104 10425 30107
rect 9180 30076 10425 30104
rect 9180 30064 9186 30076
rect 10413 30073 10425 30076
rect 10459 30073 10471 30107
rect 12360 30104 12388 30203
rect 12986 30200 12992 30252
rect 13044 30240 13050 30252
rect 13173 30243 13231 30249
rect 13173 30240 13185 30243
rect 13044 30212 13185 30240
rect 13044 30200 13050 30212
rect 13173 30209 13185 30212
rect 13219 30209 13231 30243
rect 13173 30203 13231 30209
rect 14461 30243 14519 30249
rect 14461 30209 14473 30243
rect 14507 30240 14519 30243
rect 14918 30240 14924 30252
rect 14507 30212 14924 30240
rect 14507 30209 14519 30212
rect 14461 30203 14519 30209
rect 14918 30200 14924 30212
rect 14976 30240 14982 30252
rect 15102 30240 15108 30252
rect 14976 30212 15108 30240
rect 14976 30200 14982 30212
rect 15102 30200 15108 30212
rect 15160 30200 15166 30252
rect 15473 30243 15531 30249
rect 15473 30209 15485 30243
rect 15519 30240 15531 30243
rect 15746 30240 15752 30252
rect 15519 30212 15752 30240
rect 15519 30209 15531 30212
rect 15473 30203 15531 30209
rect 15746 30200 15752 30212
rect 15804 30200 15810 30252
rect 16301 30243 16359 30249
rect 16301 30209 16313 30243
rect 16347 30240 16359 30243
rect 17034 30240 17040 30252
rect 16347 30212 17040 30240
rect 16347 30209 16359 30212
rect 16301 30203 16359 30209
rect 17034 30200 17040 30212
rect 17092 30200 17098 30252
rect 18046 30200 18052 30252
rect 18104 30240 18110 30252
rect 18233 30243 18291 30249
rect 18233 30240 18245 30243
rect 18104 30212 18245 30240
rect 18104 30200 18110 30212
rect 18233 30209 18245 30212
rect 18279 30209 18291 30243
rect 18506 30240 18512 30252
rect 18467 30212 18512 30240
rect 18233 30203 18291 30209
rect 18506 30200 18512 30212
rect 18564 30200 18570 30252
rect 19076 30249 19104 30280
rect 19337 30277 19349 30311
rect 19383 30308 19395 30311
rect 19426 30308 19432 30320
rect 19383 30280 19432 30308
rect 19383 30277 19395 30280
rect 19337 30271 19395 30277
rect 19426 30268 19432 30280
rect 19484 30268 19490 30320
rect 20346 30268 20352 30320
rect 20404 30268 20410 30320
rect 20806 30268 20812 30320
rect 20864 30308 20870 30320
rect 22112 30308 22140 30348
rect 20864 30280 22140 30308
rect 22189 30311 22247 30317
rect 20864 30268 20870 30280
rect 22189 30277 22201 30311
rect 22235 30308 22247 30311
rect 22278 30308 22284 30320
rect 22235 30280 22284 30308
rect 22235 30277 22247 30280
rect 22189 30271 22247 30277
rect 22278 30268 22284 30280
rect 22336 30268 22342 30320
rect 22388 30308 22416 30348
rect 25409 30345 25421 30379
rect 25455 30376 25467 30379
rect 25958 30376 25964 30388
rect 25455 30348 25964 30376
rect 25455 30345 25467 30348
rect 25409 30339 25467 30345
rect 25958 30336 25964 30348
rect 26016 30336 26022 30388
rect 27249 30379 27307 30385
rect 27249 30345 27261 30379
rect 27295 30376 27307 30379
rect 27338 30376 27344 30388
rect 27295 30348 27344 30376
rect 27295 30345 27307 30348
rect 27249 30339 27307 30345
rect 27338 30336 27344 30348
rect 27396 30336 27402 30388
rect 27586 30348 27936 30376
rect 27586 30308 27614 30348
rect 22388 30280 27614 30308
rect 27908 30308 27936 30348
rect 28350 30336 28356 30388
rect 28408 30376 28414 30388
rect 28408 30348 28764 30376
rect 28408 30336 28414 30348
rect 28442 30308 28448 30320
rect 27908 30280 28448 30308
rect 28442 30268 28448 30280
rect 28500 30268 28506 30320
rect 28736 30317 28764 30348
rect 28902 30336 28908 30388
rect 28960 30376 28966 30388
rect 28960 30348 29224 30376
rect 28960 30336 28966 30348
rect 28721 30311 28779 30317
rect 28721 30277 28733 30311
rect 28767 30277 28779 30311
rect 29196 30308 29224 30348
rect 29270 30336 29276 30388
rect 29328 30376 29334 30388
rect 29328 30348 29868 30376
rect 29328 30336 29334 30348
rect 29840 30317 29868 30348
rect 29609 30311 29667 30317
rect 29609 30308 29621 30311
rect 29196 30280 29621 30308
rect 28721 30271 28779 30277
rect 29609 30277 29621 30280
rect 29655 30277 29667 30311
rect 29609 30271 29667 30277
rect 29825 30311 29883 30317
rect 29825 30277 29837 30311
rect 29871 30277 29883 30311
rect 29825 30271 29883 30277
rect 19061 30243 19119 30249
rect 19061 30209 19073 30243
rect 19107 30209 19119 30243
rect 19061 30203 19119 30209
rect 21453 30243 21511 30249
rect 21453 30209 21465 30243
rect 21499 30240 21511 30243
rect 22370 30240 22376 30252
rect 21499 30212 22376 30240
rect 21499 30209 21511 30212
rect 21453 30203 21511 30209
rect 22370 30200 22376 30212
rect 22428 30200 22434 30252
rect 22465 30243 22523 30249
rect 22465 30209 22477 30243
rect 22511 30209 22523 30243
rect 23842 30240 23848 30252
rect 23803 30212 23848 30240
rect 22465 30203 22523 30209
rect 12434 30132 12440 30184
rect 12492 30172 12498 30184
rect 13449 30175 13507 30181
rect 13449 30172 13461 30175
rect 12492 30144 13461 30172
rect 12492 30132 12498 30144
rect 13449 30141 13461 30144
rect 13495 30172 13507 30175
rect 14274 30172 14280 30184
rect 13495 30144 14280 30172
rect 13495 30141 13507 30144
rect 13449 30135 13507 30141
rect 14274 30132 14280 30144
rect 14332 30132 14338 30184
rect 15562 30132 15568 30184
rect 15620 30172 15626 30184
rect 16206 30172 16212 30184
rect 15620 30144 16212 30172
rect 15620 30132 15626 30144
rect 16206 30132 16212 30144
rect 16264 30172 16270 30184
rect 17405 30175 17463 30181
rect 17405 30172 17417 30175
rect 16264 30144 17417 30172
rect 16264 30132 16270 30144
rect 17405 30141 17417 30144
rect 17451 30172 17463 30175
rect 19978 30172 19984 30184
rect 17451 30144 19984 30172
rect 17451 30141 17463 30144
rect 17405 30135 17463 30141
rect 19978 30132 19984 30144
rect 20036 30132 20042 30184
rect 20806 30172 20812 30184
rect 20767 30144 20812 30172
rect 20806 30132 20812 30144
rect 20864 30132 20870 30184
rect 22480 30172 22508 30203
rect 23842 30200 23848 30212
rect 23900 30200 23906 30252
rect 23937 30243 23995 30249
rect 23937 30209 23949 30243
rect 23983 30240 23995 30243
rect 25038 30240 25044 30252
rect 23983 30212 25044 30240
rect 23983 30209 23995 30212
rect 23937 30203 23995 30209
rect 25038 30200 25044 30212
rect 25096 30200 25102 30252
rect 26237 30243 26295 30249
rect 26237 30209 26249 30243
rect 26283 30240 26295 30243
rect 26786 30240 26792 30252
rect 26283 30212 26792 30240
rect 26283 30209 26295 30212
rect 26237 30203 26295 30209
rect 26786 30200 26792 30212
rect 26844 30200 26850 30252
rect 27246 30200 27252 30252
rect 27304 30240 27310 30252
rect 27525 30243 27583 30249
rect 27525 30240 27537 30243
rect 27304 30212 27537 30240
rect 27304 30200 27310 30212
rect 27525 30209 27537 30212
rect 27571 30209 27583 30243
rect 27525 30203 27583 30209
rect 27614 30243 27672 30249
rect 27614 30209 27626 30243
rect 27660 30209 27672 30243
rect 27614 30203 27672 30209
rect 27714 30243 27772 30249
rect 27714 30209 27726 30243
rect 27760 30209 27772 30243
rect 27714 30203 27772 30209
rect 27893 30243 27951 30249
rect 27893 30209 27905 30243
rect 27939 30240 27951 30243
rect 28166 30240 28172 30252
rect 27939 30212 28172 30240
rect 27939 30209 27951 30212
rect 27893 30203 27951 30209
rect 23750 30172 23756 30184
rect 22066 30144 23756 30172
rect 22066 30104 22094 30144
rect 23750 30132 23756 30144
rect 23808 30132 23814 30184
rect 24026 30172 24032 30184
rect 23987 30144 24032 30172
rect 24026 30132 24032 30144
rect 24084 30132 24090 30184
rect 24854 30172 24860 30184
rect 24815 30144 24860 30172
rect 24854 30132 24860 30144
rect 24912 30132 24918 30184
rect 24949 30175 25007 30181
rect 24949 30141 24961 30175
rect 24995 30141 25007 30175
rect 24949 30135 25007 30141
rect 12360 30076 17264 30104
rect 10413 30067 10471 30073
rect 9953 30039 10011 30045
rect 9953 30005 9965 30039
rect 9999 30036 10011 30039
rect 10134 30036 10140 30048
rect 9999 30008 10140 30036
rect 9999 30005 10011 30008
rect 9953 29999 10011 30005
rect 10134 29996 10140 30008
rect 10192 29996 10198 30048
rect 11606 29996 11612 30048
rect 11664 30036 11670 30048
rect 12805 30039 12863 30045
rect 12805 30036 12817 30039
rect 11664 30008 12817 30036
rect 11664 29996 11670 30008
rect 12805 30005 12817 30008
rect 12851 30005 12863 30039
rect 15286 30036 15292 30048
rect 15247 30008 15292 30036
rect 12805 29999 12863 30005
rect 15286 29996 15292 30008
rect 15344 29996 15350 30048
rect 16850 30036 16856 30048
rect 16811 30008 16856 30036
rect 16850 29996 16856 30008
rect 16908 29996 16914 30048
rect 17236 30036 17264 30076
rect 20364 30076 22094 30104
rect 20364 30036 20392 30076
rect 23566 30064 23572 30116
rect 23624 30104 23630 30116
rect 24964 30104 24992 30135
rect 27629 30116 27657 30203
rect 23624 30076 24992 30104
rect 23624 30064 23630 30076
rect 27614 30064 27620 30116
rect 27672 30064 27678 30116
rect 17236 30008 20392 30036
rect 21174 29996 21180 30048
rect 21232 30036 21238 30048
rect 21269 30039 21327 30045
rect 21269 30036 21281 30039
rect 21232 30008 21281 30036
rect 21232 29996 21238 30008
rect 21269 30005 21281 30008
rect 21315 30005 21327 30039
rect 23474 30036 23480 30048
rect 23435 30008 23480 30036
rect 21269 29999 21327 30005
rect 23474 29996 23480 30008
rect 23532 29996 23538 30048
rect 24854 29996 24860 30048
rect 24912 30036 24918 30048
rect 25961 30039 26019 30045
rect 25961 30036 25973 30039
rect 24912 30008 25973 30036
rect 24912 29996 24918 30008
rect 25961 30005 25973 30008
rect 26007 30005 26019 30039
rect 27724 30036 27752 30203
rect 28166 30200 28172 30212
rect 28224 30200 28230 30252
rect 28534 30249 28540 30252
rect 28532 30240 28540 30249
rect 28495 30212 28540 30240
rect 28532 30203 28540 30212
rect 28534 30200 28540 30203
rect 28592 30200 28598 30252
rect 28626 30200 28632 30252
rect 28684 30240 28690 30252
rect 28684 30212 28729 30240
rect 28684 30200 28690 30212
rect 28810 30200 28816 30252
rect 28868 30249 28874 30252
rect 28868 30243 28907 30249
rect 28895 30209 28907 30243
rect 28997 30243 29055 30249
rect 28997 30240 29009 30243
rect 28868 30203 28907 30209
rect 28940 30212 29009 30240
rect 28868 30200 28874 30203
rect 28940 30116 28968 30212
rect 28997 30209 29009 30212
rect 29043 30209 29055 30243
rect 28997 30203 29055 30209
rect 30653 30243 30711 30249
rect 30653 30209 30665 30243
rect 30699 30240 30711 30243
rect 30926 30240 30932 30252
rect 30699 30212 30932 30240
rect 30699 30209 30711 30212
rect 30653 30203 30711 30209
rect 30926 30200 30932 30212
rect 30984 30200 30990 30252
rect 31478 30240 31484 30252
rect 31439 30212 31484 30240
rect 31478 30200 31484 30212
rect 31536 30200 31542 30252
rect 32122 30200 32128 30252
rect 32180 30240 32186 30252
rect 32309 30243 32367 30249
rect 32309 30240 32321 30243
rect 32180 30212 32321 30240
rect 32180 30200 32186 30212
rect 32309 30209 32321 30212
rect 32355 30209 32367 30243
rect 32309 30203 32367 30209
rect 33042 30200 33048 30252
rect 33100 30240 33106 30252
rect 33669 30243 33727 30249
rect 33669 30240 33681 30243
rect 33100 30212 33681 30240
rect 33100 30200 33106 30212
rect 33669 30209 33681 30212
rect 33715 30209 33727 30243
rect 33669 30203 33727 30209
rect 33962 30200 33968 30252
rect 34020 30240 34026 30252
rect 34020 30212 34468 30240
rect 34020 30200 34026 30212
rect 30558 30172 30564 30184
rect 30519 30144 30564 30172
rect 30558 30132 30564 30144
rect 30616 30132 30622 30184
rect 31021 30175 31079 30181
rect 31021 30141 31033 30175
rect 31067 30172 31079 30175
rect 31570 30172 31576 30184
rect 31067 30144 31576 30172
rect 31067 30141 31079 30144
rect 31021 30135 31079 30141
rect 31570 30132 31576 30144
rect 31628 30132 31634 30184
rect 32585 30175 32643 30181
rect 32585 30141 32597 30175
rect 32631 30172 32643 30175
rect 33318 30172 33324 30184
rect 32631 30144 33324 30172
rect 32631 30141 32643 30144
rect 32585 30135 32643 30141
rect 33318 30132 33324 30144
rect 33376 30132 33382 30184
rect 33413 30175 33471 30181
rect 33413 30141 33425 30175
rect 33459 30141 33471 30175
rect 33413 30135 33471 30141
rect 27890 30064 27896 30116
rect 27948 30104 27954 30116
rect 27948 30076 28488 30104
rect 27948 30064 27954 30076
rect 28074 30036 28080 30048
rect 27724 30008 28080 30036
rect 25961 29999 26019 30005
rect 28074 29996 28080 30008
rect 28132 29996 28138 30048
rect 28350 30036 28356 30048
rect 28311 30008 28356 30036
rect 28350 29996 28356 30008
rect 28408 29996 28414 30048
rect 28460 30036 28488 30076
rect 28902 30064 28908 30116
rect 28960 30076 28968 30116
rect 28960 30064 28966 30076
rect 29086 30064 29092 30116
rect 29144 30104 29150 30116
rect 29457 30107 29515 30113
rect 29457 30104 29469 30107
rect 29144 30076 29469 30104
rect 29144 30064 29150 30076
rect 29457 30073 29469 30076
rect 29503 30073 29515 30107
rect 29457 30067 29515 30073
rect 29564 30076 31616 30104
rect 29564 30036 29592 30076
rect 28460 30008 29592 30036
rect 29641 30039 29699 30045
rect 29641 30005 29653 30039
rect 29687 30036 29699 30039
rect 29730 30036 29736 30048
rect 29687 30008 29736 30036
rect 29687 30005 29699 30008
rect 29641 29999 29699 30005
rect 29730 29996 29736 30008
rect 29788 29996 29794 30048
rect 31588 30045 31616 30076
rect 31573 30039 31631 30045
rect 31573 30005 31585 30039
rect 31619 30005 31631 30039
rect 33428 30036 33456 30135
rect 34440 30104 34468 30212
rect 34793 30107 34851 30113
rect 34793 30104 34805 30107
rect 34440 30076 34805 30104
rect 34793 30073 34805 30076
rect 34839 30073 34851 30107
rect 34793 30067 34851 30073
rect 34422 30036 34428 30048
rect 33428 30008 34428 30036
rect 31573 29999 31631 30005
rect 34422 29996 34428 30008
rect 34480 29996 34486 30048
rect 1104 29946 37628 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 37628 29946
rect 1104 29872 37628 29894
rect 6914 29792 6920 29844
rect 6972 29832 6978 29844
rect 6972 29804 8616 29832
rect 6972 29792 6978 29804
rect 7837 29767 7895 29773
rect 7837 29764 7849 29767
rect 6886 29736 7849 29764
rect 6886 29696 6914 29736
rect 7837 29733 7849 29736
rect 7883 29733 7895 29767
rect 7837 29727 7895 29733
rect 8018 29724 8024 29776
rect 8076 29764 8082 29776
rect 8076 29736 8432 29764
rect 8076 29724 8082 29736
rect 8294 29696 8300 29708
rect 5920 29668 6914 29696
rect 8255 29668 8300 29696
rect 5920 29637 5948 29668
rect 8294 29656 8300 29668
rect 8352 29656 8358 29708
rect 8404 29705 8432 29736
rect 8389 29699 8447 29705
rect 8389 29665 8401 29699
rect 8435 29665 8447 29699
rect 8389 29659 8447 29665
rect 5905 29631 5963 29637
rect 5905 29597 5917 29631
rect 5951 29597 5963 29631
rect 5905 29591 5963 29597
rect 6549 29631 6607 29637
rect 6549 29597 6561 29631
rect 6595 29628 6607 29631
rect 6914 29628 6920 29640
rect 6595 29600 6920 29628
rect 6595 29597 6607 29600
rect 6549 29591 6607 29597
rect 6914 29588 6920 29600
rect 6972 29588 6978 29640
rect 7193 29631 7251 29637
rect 7193 29597 7205 29631
rect 7239 29628 7251 29631
rect 8588 29628 8616 29804
rect 8754 29792 8760 29844
rect 8812 29832 8818 29844
rect 9214 29832 9220 29844
rect 8812 29804 9220 29832
rect 8812 29792 8818 29804
rect 9214 29792 9220 29804
rect 9272 29832 9278 29844
rect 12894 29832 12900 29844
rect 9272 29804 12756 29832
rect 12855 29804 12900 29832
rect 9272 29792 9278 29804
rect 11146 29764 11152 29776
rect 10244 29736 11152 29764
rect 10244 29705 10272 29736
rect 11146 29724 11152 29736
rect 11204 29724 11210 29776
rect 10229 29699 10287 29705
rect 10229 29665 10241 29699
rect 10275 29665 10287 29699
rect 10229 29659 10287 29665
rect 10413 29699 10471 29705
rect 10413 29665 10425 29699
rect 10459 29696 10471 29699
rect 10870 29696 10876 29708
rect 10459 29668 10876 29696
rect 10459 29665 10471 29668
rect 10413 29659 10471 29665
rect 10870 29656 10876 29668
rect 10928 29656 10934 29708
rect 11054 29656 11060 29708
rect 11112 29696 11118 29708
rect 11425 29699 11483 29705
rect 11425 29696 11437 29699
rect 11112 29668 11437 29696
rect 11112 29656 11118 29668
rect 11425 29665 11437 29668
rect 11471 29665 11483 29699
rect 12728 29696 12756 29804
rect 12894 29792 12900 29804
rect 12952 29792 12958 29844
rect 14553 29835 14611 29841
rect 14553 29801 14565 29835
rect 14599 29832 14611 29835
rect 15562 29832 15568 29844
rect 14599 29804 15568 29832
rect 14599 29801 14611 29804
rect 14553 29795 14611 29801
rect 15562 29792 15568 29804
rect 15620 29792 15626 29844
rect 15746 29832 15752 29844
rect 15707 29804 15752 29832
rect 15746 29792 15752 29804
rect 15804 29792 15810 29844
rect 19702 29832 19708 29844
rect 18340 29804 19564 29832
rect 19663 29804 19708 29832
rect 13630 29724 13636 29776
rect 13688 29764 13694 29776
rect 18340 29764 18368 29804
rect 13688 29736 18368 29764
rect 19536 29764 19564 29804
rect 19702 29792 19708 29804
rect 19760 29792 19766 29844
rect 22278 29832 22284 29844
rect 19812 29804 22284 29832
rect 19812 29764 19840 29804
rect 22278 29792 22284 29804
rect 22336 29792 22342 29844
rect 22370 29792 22376 29844
rect 22428 29832 22434 29844
rect 23109 29835 23167 29841
rect 23109 29832 23121 29835
rect 22428 29804 23121 29832
rect 22428 29792 22434 29804
rect 23109 29801 23121 29804
rect 23155 29801 23167 29835
rect 23109 29795 23167 29801
rect 25038 29792 25044 29844
rect 25096 29832 25102 29844
rect 26697 29835 26755 29841
rect 26697 29832 26709 29835
rect 25096 29804 26709 29832
rect 25096 29792 25102 29804
rect 26697 29801 26709 29804
rect 26743 29832 26755 29835
rect 27430 29832 27436 29844
rect 26743 29804 27436 29832
rect 26743 29801 26755 29804
rect 26697 29795 26755 29801
rect 27430 29792 27436 29804
rect 27488 29792 27494 29844
rect 28445 29835 28503 29841
rect 28445 29801 28457 29835
rect 28491 29832 28503 29835
rect 28902 29832 28908 29844
rect 28491 29804 28908 29832
rect 28491 29801 28503 29804
rect 28445 29795 28503 29801
rect 28902 29792 28908 29804
rect 28960 29792 28966 29844
rect 30929 29835 30987 29841
rect 30929 29832 30941 29835
rect 30116 29804 30941 29832
rect 19536 29736 19840 29764
rect 13688 29724 13694 29736
rect 16393 29699 16451 29705
rect 12728 29668 13768 29696
rect 11425 29659 11483 29665
rect 9125 29631 9183 29637
rect 9125 29628 9137 29631
rect 7239 29600 8524 29628
rect 8588 29600 9137 29628
rect 7239 29597 7251 29600
rect 7193 29591 7251 29597
rect 6086 29492 6092 29504
rect 6047 29464 6092 29492
rect 6086 29452 6092 29464
rect 6144 29452 6150 29504
rect 6641 29495 6699 29501
rect 6641 29461 6653 29495
rect 6687 29492 6699 29495
rect 7282 29492 7288 29504
rect 6687 29464 7288 29492
rect 6687 29461 6699 29464
rect 6641 29455 6699 29461
rect 7282 29452 7288 29464
rect 7340 29452 7346 29504
rect 7377 29495 7435 29501
rect 7377 29461 7389 29495
rect 7423 29492 7435 29495
rect 8110 29492 8116 29504
rect 7423 29464 8116 29492
rect 7423 29461 7435 29464
rect 7377 29455 7435 29461
rect 8110 29452 8116 29464
rect 8168 29452 8174 29504
rect 8205 29495 8263 29501
rect 8205 29461 8217 29495
rect 8251 29492 8263 29495
rect 8386 29492 8392 29504
rect 8251 29464 8392 29492
rect 8251 29461 8263 29464
rect 8205 29455 8263 29461
rect 8386 29452 8392 29464
rect 8444 29452 8450 29504
rect 8496 29492 8524 29600
rect 9125 29597 9137 29600
rect 9171 29597 9183 29631
rect 10134 29628 10140 29640
rect 10095 29600 10140 29628
rect 9125 29591 9183 29597
rect 10134 29588 10140 29600
rect 10192 29588 10198 29640
rect 11146 29628 11152 29640
rect 11107 29600 11152 29628
rect 11146 29588 11152 29600
rect 11204 29588 11210 29640
rect 13740 29637 13768 29668
rect 16393 29665 16405 29699
rect 16439 29696 16451 29699
rect 18138 29696 18144 29708
rect 16439 29668 18144 29696
rect 16439 29665 16451 29668
rect 16393 29659 16451 29665
rect 18138 29656 18144 29668
rect 18196 29696 18202 29708
rect 18233 29699 18291 29705
rect 18233 29696 18245 29699
rect 18196 29668 18245 29696
rect 18196 29656 18202 29668
rect 18233 29665 18245 29668
rect 18279 29665 18291 29699
rect 18233 29659 18291 29665
rect 13725 29631 13783 29637
rect 13725 29597 13737 29631
rect 13771 29628 13783 29631
rect 17037 29631 17095 29637
rect 13771 29600 15516 29628
rect 13771 29597 13783 29600
rect 13725 29591 13783 29597
rect 15488 29572 15516 29600
rect 17037 29597 17049 29631
rect 17083 29628 17095 29631
rect 17494 29628 17500 29640
rect 17083 29600 17500 29628
rect 17083 29597 17095 29600
rect 17037 29591 17095 29597
rect 17494 29588 17500 29600
rect 17552 29628 17558 29640
rect 18506 29628 18512 29640
rect 17552 29600 18512 29628
rect 17552 29588 17558 29600
rect 18506 29588 18512 29600
rect 18564 29588 18570 29640
rect 18598 29588 18604 29640
rect 18656 29628 18662 29640
rect 19812 29637 19840 29736
rect 22649 29767 22707 29773
rect 22649 29733 22661 29767
rect 22695 29764 22707 29767
rect 22695 29736 23612 29764
rect 22695 29733 22707 29736
rect 22649 29727 22707 29733
rect 23584 29708 23612 29736
rect 27706 29724 27712 29776
rect 27764 29764 27770 29776
rect 27764 29736 28120 29764
rect 27764 29724 27770 29736
rect 20901 29699 20959 29705
rect 20901 29665 20913 29699
rect 20947 29696 20959 29699
rect 22922 29696 22928 29708
rect 20947 29668 22928 29696
rect 20947 29665 20959 29668
rect 20901 29659 20959 29665
rect 22922 29656 22928 29668
rect 22980 29656 22986 29708
rect 23566 29696 23572 29708
rect 23527 29668 23572 29696
rect 23566 29656 23572 29668
rect 23624 29656 23630 29708
rect 23658 29656 23664 29708
rect 23716 29696 23722 29708
rect 25222 29696 25228 29708
rect 23716 29668 23761 29696
rect 25183 29668 25228 29696
rect 23716 29656 23722 29668
rect 25222 29656 25228 29668
rect 25280 29656 25286 29708
rect 27982 29696 27988 29708
rect 27943 29668 27988 29696
rect 27982 29656 27988 29668
rect 28040 29656 28046 29708
rect 28092 29705 28120 29736
rect 28258 29724 28264 29776
rect 28316 29764 28322 29776
rect 29914 29764 29920 29776
rect 28316 29736 29920 29764
rect 28316 29724 28322 29736
rect 29914 29724 29920 29736
rect 29972 29764 29978 29776
rect 30116 29764 30144 29804
rect 30929 29801 30941 29804
rect 30975 29801 30987 29835
rect 33042 29832 33048 29844
rect 33003 29804 33048 29832
rect 30929 29795 30987 29801
rect 33042 29792 33048 29804
rect 33100 29792 33106 29844
rect 29972 29736 30144 29764
rect 29972 29724 29978 29736
rect 28077 29699 28135 29705
rect 28077 29665 28089 29699
rect 28123 29696 28135 29699
rect 28442 29696 28448 29708
rect 28123 29668 28448 29696
rect 28123 29665 28135 29668
rect 28077 29659 28135 29665
rect 28442 29656 28448 29668
rect 28500 29656 28506 29708
rect 28905 29699 28963 29705
rect 28905 29665 28917 29699
rect 28951 29696 28963 29699
rect 28994 29696 29000 29708
rect 28951 29668 29000 29696
rect 28951 29665 28963 29668
rect 28905 29659 28963 29665
rect 28994 29656 29000 29668
rect 29052 29656 29058 29708
rect 33873 29699 33931 29705
rect 33873 29665 33885 29699
rect 33919 29696 33931 29699
rect 33962 29696 33968 29708
rect 33919 29668 33968 29696
rect 33919 29665 33931 29668
rect 33873 29659 33931 29665
rect 33962 29656 33968 29668
rect 34020 29656 34026 29708
rect 19797 29631 19855 29637
rect 18656 29600 19748 29628
rect 18656 29588 18662 29600
rect 9217 29563 9275 29569
rect 9217 29529 9229 29563
rect 9263 29560 9275 29563
rect 14642 29560 14648 29572
rect 9263 29532 10548 29560
rect 9263 29529 9275 29532
rect 9217 29523 9275 29529
rect 9769 29495 9827 29501
rect 9769 29492 9781 29495
rect 8496 29464 9781 29492
rect 9769 29461 9781 29464
rect 9815 29461 9827 29495
rect 10520 29492 10548 29532
rect 11532 29532 11914 29560
rect 14603 29532 14648 29560
rect 11532 29492 11560 29532
rect 14642 29520 14648 29532
rect 14700 29520 14706 29572
rect 15470 29520 15476 29572
rect 15528 29560 15534 29572
rect 17313 29563 17371 29569
rect 17313 29560 17325 29563
rect 15528 29532 17325 29560
rect 15528 29520 15534 29532
rect 17313 29529 17325 29532
rect 17359 29560 17371 29563
rect 19610 29560 19616 29572
rect 17359 29532 19616 29560
rect 17359 29529 17371 29532
rect 17313 29523 17371 29529
rect 19610 29520 19616 29532
rect 19668 29520 19674 29572
rect 19720 29560 19748 29600
rect 19797 29597 19809 29631
rect 19843 29597 19855 29631
rect 23474 29628 23480 29640
rect 23435 29600 23480 29628
rect 19797 29591 19855 29597
rect 23474 29588 23480 29600
rect 23532 29588 23538 29640
rect 24854 29588 24860 29640
rect 24912 29628 24918 29640
rect 24949 29631 25007 29637
rect 24949 29628 24961 29631
rect 24912 29600 24961 29628
rect 24912 29588 24918 29600
rect 24949 29597 24961 29600
rect 24995 29597 25007 29631
rect 24949 29591 25007 29597
rect 27709 29631 27767 29637
rect 27709 29597 27721 29631
rect 27755 29628 27767 29631
rect 27798 29628 27804 29640
rect 27755 29600 27804 29628
rect 27755 29597 27767 29600
rect 27709 29591 27767 29597
rect 27798 29588 27804 29600
rect 27856 29588 27862 29640
rect 27890 29588 27896 29640
rect 27948 29628 27954 29640
rect 28261 29631 28319 29637
rect 27948 29600 27993 29628
rect 27948 29588 27954 29600
rect 28261 29597 28273 29631
rect 28307 29628 28319 29631
rect 28810 29628 28816 29640
rect 28307 29600 28816 29628
rect 28307 29597 28319 29600
rect 28261 29591 28319 29597
rect 21174 29560 21180 29572
rect 19720 29532 20392 29560
rect 21135 29532 21180 29560
rect 13630 29492 13636 29504
rect 10520 29464 11560 29492
rect 13591 29464 13636 29492
rect 9769 29455 9827 29461
rect 13630 29452 13636 29464
rect 13688 29452 13694 29504
rect 16114 29492 16120 29504
rect 16075 29464 16120 29492
rect 16114 29452 16120 29464
rect 16172 29452 16178 29504
rect 16209 29495 16267 29501
rect 16209 29461 16221 29495
rect 16255 29492 16267 29495
rect 16298 29492 16304 29504
rect 16255 29464 16304 29492
rect 16255 29461 16267 29464
rect 16209 29455 16267 29461
rect 16298 29452 16304 29464
rect 16356 29452 16362 29504
rect 18414 29492 18420 29504
rect 18375 29464 18420 29492
rect 18414 29452 18420 29464
rect 18472 29452 18478 29504
rect 18506 29452 18512 29504
rect 18564 29492 18570 29504
rect 18877 29495 18935 29501
rect 18564 29464 18609 29492
rect 18564 29452 18570 29464
rect 18877 29461 18889 29495
rect 18923 29492 18935 29495
rect 20254 29492 20260 29504
rect 18923 29464 20260 29492
rect 18923 29461 18935 29464
rect 18877 29455 18935 29461
rect 20254 29452 20260 29464
rect 20312 29452 20318 29504
rect 20364 29492 20392 29532
rect 21174 29520 21180 29532
rect 21232 29520 21238 29572
rect 21634 29520 21640 29572
rect 21692 29520 21698 29572
rect 26510 29560 26516 29572
rect 26450 29532 26516 29560
rect 26510 29520 26516 29532
rect 26568 29520 26574 29572
rect 28074 29520 28080 29572
rect 28132 29560 28138 29572
rect 28276 29560 28304 29591
rect 28810 29588 28816 29600
rect 28868 29588 28874 29640
rect 29086 29628 29092 29640
rect 29047 29600 29092 29628
rect 29086 29588 29092 29600
rect 29144 29588 29150 29640
rect 29178 29588 29184 29640
rect 29236 29628 29242 29640
rect 29236 29600 29281 29628
rect 29236 29588 29242 29600
rect 29546 29588 29552 29640
rect 29604 29628 29610 29640
rect 29733 29631 29791 29637
rect 29733 29628 29745 29631
rect 29604 29600 29745 29628
rect 29604 29588 29610 29600
rect 29733 29597 29745 29600
rect 29779 29597 29791 29631
rect 29733 29591 29791 29597
rect 29822 29588 29828 29640
rect 29880 29628 29886 29640
rect 30101 29631 30159 29637
rect 30101 29628 30113 29631
rect 29880 29600 30113 29628
rect 29880 29588 29886 29600
rect 30101 29597 30113 29600
rect 30147 29597 30159 29631
rect 30101 29591 30159 29597
rect 31757 29631 31815 29637
rect 31757 29597 31769 29631
rect 31803 29628 31815 29631
rect 32030 29628 32036 29640
rect 31803 29600 32036 29628
rect 31803 29597 31815 29600
rect 31757 29591 31815 29597
rect 32030 29588 32036 29600
rect 32088 29588 32094 29640
rect 32214 29628 32220 29640
rect 32175 29600 32220 29628
rect 32214 29588 32220 29600
rect 32272 29588 32278 29640
rect 32861 29631 32919 29637
rect 32861 29597 32873 29631
rect 32907 29628 32919 29631
rect 33505 29631 33563 29637
rect 33505 29628 33517 29631
rect 32907 29600 33517 29628
rect 32907 29597 32919 29600
rect 32861 29591 32919 29597
rect 33505 29597 33517 29600
rect 33551 29597 33563 29631
rect 33505 29591 33563 29597
rect 33689 29631 33747 29637
rect 33689 29597 33701 29631
rect 33735 29597 33747 29631
rect 33689 29591 33747 29597
rect 28132 29532 28304 29560
rect 28905 29563 28963 29569
rect 28132 29520 28138 29532
rect 28905 29529 28917 29563
rect 28951 29560 28963 29563
rect 29917 29563 29975 29569
rect 29917 29560 29929 29563
rect 28951 29532 29929 29560
rect 28951 29529 28963 29532
rect 28905 29523 28963 29529
rect 29917 29529 29929 29532
rect 29963 29529 29975 29563
rect 29917 29523 29975 29529
rect 30006 29520 30012 29572
rect 30064 29560 30070 29572
rect 30742 29560 30748 29572
rect 30064 29532 30109 29560
rect 30703 29532 30748 29560
rect 30064 29520 30070 29532
rect 30742 29520 30748 29532
rect 30800 29520 30806 29572
rect 31665 29563 31723 29569
rect 31665 29529 31677 29563
rect 31711 29560 31723 29563
rect 33410 29560 33416 29572
rect 31711 29532 33416 29560
rect 31711 29529 31723 29532
rect 31665 29523 31723 29529
rect 33410 29520 33416 29532
rect 33468 29520 33474 29572
rect 26786 29492 26792 29504
rect 20364 29464 26792 29492
rect 26786 29452 26792 29464
rect 26844 29452 26850 29504
rect 29730 29452 29736 29504
rect 29788 29492 29794 29504
rect 30285 29495 30343 29501
rect 30285 29492 30297 29495
rect 29788 29464 30297 29492
rect 29788 29452 29794 29464
rect 30285 29461 30297 29464
rect 30331 29461 30343 29495
rect 30285 29455 30343 29461
rect 30650 29452 30656 29504
rect 30708 29492 30714 29504
rect 30945 29495 31003 29501
rect 30945 29492 30957 29495
rect 30708 29464 30957 29492
rect 30708 29452 30714 29464
rect 30945 29461 30957 29464
rect 30991 29461 31003 29495
rect 31110 29492 31116 29504
rect 31071 29464 31116 29492
rect 30945 29455 31003 29461
rect 31110 29452 31116 29464
rect 31168 29452 31174 29504
rect 32398 29492 32404 29504
rect 32359 29464 32404 29492
rect 32398 29452 32404 29464
rect 32456 29452 32462 29504
rect 33226 29452 33232 29504
rect 33284 29492 33290 29504
rect 33704 29492 33732 29591
rect 33284 29464 33732 29492
rect 33284 29452 33290 29464
rect 1104 29402 37628 29424
rect 1104 29350 4874 29402
rect 4926 29350 4938 29402
rect 4990 29350 5002 29402
rect 5054 29350 5066 29402
rect 5118 29350 5130 29402
rect 5182 29350 35594 29402
rect 35646 29350 35658 29402
rect 35710 29350 35722 29402
rect 35774 29350 35786 29402
rect 35838 29350 35850 29402
rect 35902 29350 37628 29402
rect 1104 29328 37628 29350
rect 9306 29248 9312 29300
rect 9364 29288 9370 29300
rect 11057 29291 11115 29297
rect 9364 29260 9996 29288
rect 9364 29248 9370 29260
rect 6086 29180 6092 29232
rect 6144 29220 6150 29232
rect 6825 29223 6883 29229
rect 6825 29220 6837 29223
rect 6144 29192 6837 29220
rect 6144 29180 6150 29192
rect 6825 29189 6837 29192
rect 6871 29189 6883 29223
rect 6825 29183 6883 29189
rect 7282 29180 7288 29232
rect 7340 29180 7346 29232
rect 8110 29180 8116 29232
rect 8168 29220 8174 29232
rect 9585 29223 9643 29229
rect 9585 29220 9597 29223
rect 8168 29192 9597 29220
rect 8168 29180 8174 29192
rect 9585 29189 9597 29192
rect 9631 29189 9643 29223
rect 9968 29220 9996 29260
rect 11057 29257 11069 29291
rect 11103 29288 11115 29291
rect 11238 29288 11244 29300
rect 11103 29260 11244 29288
rect 11103 29257 11115 29260
rect 11057 29251 11115 29257
rect 11238 29248 11244 29260
rect 11296 29248 11302 29300
rect 14642 29248 14648 29300
rect 14700 29288 14706 29300
rect 17221 29291 17279 29297
rect 14700 29260 16160 29288
rect 14700 29248 14706 29260
rect 9968 29192 10074 29220
rect 9585 29183 9643 29189
rect 13630 29180 13636 29232
rect 13688 29180 13694 29232
rect 15562 29180 15568 29232
rect 15620 29180 15626 29232
rect 6454 29112 6460 29164
rect 6512 29152 6518 29164
rect 6549 29155 6607 29161
rect 6549 29152 6561 29155
rect 6512 29124 6561 29152
rect 6512 29112 6518 29124
rect 6549 29121 6561 29124
rect 6595 29121 6607 29155
rect 6549 29115 6607 29121
rect 11698 29112 11704 29164
rect 11756 29152 11762 29164
rect 11885 29155 11943 29161
rect 11885 29152 11897 29155
rect 11756 29124 11897 29152
rect 11756 29112 11762 29124
rect 11885 29121 11897 29124
rect 11931 29121 11943 29155
rect 11885 29115 11943 29121
rect 9306 29084 9312 29096
rect 9267 29056 9312 29084
rect 9306 29044 9312 29056
rect 9364 29044 9370 29096
rect 11146 29044 11152 29096
rect 11204 29084 11210 29096
rect 12345 29087 12403 29093
rect 12345 29084 12357 29087
rect 11204 29056 12357 29084
rect 11204 29044 11210 29056
rect 12345 29053 12357 29056
rect 12391 29053 12403 29087
rect 12618 29084 12624 29096
rect 12579 29056 12624 29084
rect 12345 29047 12403 29053
rect 11790 29016 11796 29028
rect 11751 28988 11796 29016
rect 11790 28976 11796 28988
rect 11848 28976 11854 29028
rect 12360 29016 12388 29047
rect 12618 29044 12624 29056
rect 12676 29044 12682 29096
rect 14550 29084 14556 29096
rect 14511 29056 14556 29084
rect 14550 29044 14556 29056
rect 14608 29044 14614 29096
rect 14829 29087 14887 29093
rect 14829 29053 14841 29087
rect 14875 29084 14887 29087
rect 15286 29084 15292 29096
rect 14875 29056 15292 29084
rect 14875 29053 14887 29056
rect 14829 29047 14887 29053
rect 15286 29044 15292 29056
rect 15344 29044 15350 29096
rect 16132 29084 16160 29260
rect 17221 29257 17233 29291
rect 17267 29288 17279 29291
rect 18414 29288 18420 29300
rect 17267 29260 18420 29288
rect 17267 29257 17279 29260
rect 17221 29251 17279 29257
rect 18414 29248 18420 29260
rect 18472 29248 18478 29300
rect 21361 29291 21419 29297
rect 21361 29257 21373 29291
rect 21407 29288 21419 29291
rect 21634 29288 21640 29300
rect 21407 29260 21640 29288
rect 21407 29257 21419 29260
rect 21361 29251 21419 29257
rect 21634 29248 21640 29260
rect 21692 29248 21698 29300
rect 22741 29291 22799 29297
rect 22741 29257 22753 29291
rect 22787 29288 22799 29291
rect 23569 29291 23627 29297
rect 23569 29288 23581 29291
rect 22787 29260 23581 29288
rect 22787 29257 22799 29260
rect 22741 29251 22799 29257
rect 23569 29257 23581 29260
rect 23615 29257 23627 29291
rect 23569 29251 23627 29257
rect 23750 29248 23756 29300
rect 23808 29288 23814 29300
rect 26694 29288 26700 29300
rect 23808 29260 26700 29288
rect 23808 29248 23814 29260
rect 26694 29248 26700 29260
rect 26752 29248 26758 29300
rect 29089 29291 29147 29297
rect 29089 29257 29101 29291
rect 29135 29288 29147 29291
rect 29178 29288 29184 29300
rect 29135 29260 29184 29288
rect 29135 29257 29147 29260
rect 29089 29251 29147 29257
rect 29178 29248 29184 29260
rect 29236 29248 29242 29300
rect 29546 29288 29552 29300
rect 29507 29260 29552 29288
rect 29546 29248 29552 29260
rect 29604 29248 29610 29300
rect 29638 29248 29644 29300
rect 29696 29288 29702 29300
rect 29733 29291 29791 29297
rect 29733 29288 29745 29291
rect 29696 29260 29745 29288
rect 29696 29248 29702 29260
rect 29733 29257 29745 29260
rect 29779 29257 29791 29291
rect 31294 29288 31300 29300
rect 31207 29260 31300 29288
rect 29733 29251 29791 29257
rect 31294 29248 31300 29260
rect 31352 29288 31358 29300
rect 31662 29288 31668 29300
rect 31352 29260 31668 29288
rect 31352 29248 31358 29260
rect 31662 29248 31668 29260
rect 31720 29248 31726 29300
rect 31757 29291 31815 29297
rect 31757 29257 31769 29291
rect 31803 29288 31815 29291
rect 32214 29288 32220 29300
rect 31803 29260 32220 29288
rect 31803 29257 31815 29260
rect 31757 29251 31815 29257
rect 32214 29248 32220 29260
rect 32272 29248 32278 29300
rect 33045 29291 33103 29297
rect 33045 29257 33057 29291
rect 33091 29288 33103 29291
rect 33134 29288 33140 29300
rect 33091 29260 33140 29288
rect 33091 29257 33103 29260
rect 33045 29251 33103 29257
rect 33134 29248 33140 29260
rect 33192 29248 33198 29300
rect 34885 29291 34943 29297
rect 34885 29257 34897 29291
rect 34931 29257 34943 29291
rect 34885 29251 34943 29257
rect 19521 29223 19579 29229
rect 19521 29220 19533 29223
rect 18262 29192 19533 29220
rect 19521 29189 19533 29192
rect 19567 29189 19579 29223
rect 26510 29220 26516 29232
rect 26358 29192 26516 29220
rect 19521 29183 19579 29189
rect 26510 29180 26516 29192
rect 26568 29180 26574 29232
rect 27525 29223 27583 29229
rect 27525 29189 27537 29223
rect 27571 29220 27583 29223
rect 30006 29220 30012 29232
rect 27571 29192 30012 29220
rect 27571 29189 27583 29192
rect 27525 29183 27583 29189
rect 30006 29180 30012 29192
rect 30064 29220 30070 29232
rect 31389 29223 31447 29229
rect 30064 29192 30236 29220
rect 30064 29180 30070 29192
rect 19610 29152 19616 29164
rect 19523 29124 19616 29152
rect 19610 29112 19616 29124
rect 19668 29112 19674 29164
rect 20254 29152 20260 29164
rect 20215 29124 20260 29152
rect 20254 29112 20260 29124
rect 20312 29112 20318 29164
rect 21453 29155 21511 29161
rect 21453 29121 21465 29155
rect 21499 29152 21511 29155
rect 22186 29152 22192 29164
rect 21499 29124 22192 29152
rect 21499 29121 21511 29124
rect 21453 29115 21511 29121
rect 22186 29112 22192 29124
rect 22244 29112 22250 29164
rect 23566 29112 23572 29164
rect 23624 29152 23630 29164
rect 23937 29155 23995 29161
rect 23937 29152 23949 29155
rect 23624 29124 23949 29152
rect 23624 29112 23630 29124
rect 23937 29121 23949 29124
rect 23983 29121 23995 29155
rect 27430 29152 27436 29164
rect 27391 29124 27436 29152
rect 23937 29115 23995 29121
rect 27430 29112 27436 29124
rect 27488 29112 27494 29164
rect 28350 29152 28356 29164
rect 28311 29124 28356 29152
rect 28350 29112 28356 29124
rect 28408 29112 28414 29164
rect 28534 29152 28540 29164
rect 28495 29124 28540 29152
rect 28534 29112 28540 29124
rect 28592 29112 28598 29164
rect 28902 29152 28908 29164
rect 28863 29124 28908 29152
rect 28902 29112 28908 29124
rect 28960 29112 28966 29164
rect 29674 29155 29732 29161
rect 29674 29152 29686 29155
rect 29012 29124 29686 29152
rect 18598 29084 18604 29096
rect 16132 29056 18604 29084
rect 18598 29044 18604 29056
rect 18656 29044 18662 29096
rect 18966 29084 18972 29096
rect 18927 29056 18972 29084
rect 18966 29044 18972 29056
rect 19024 29044 19030 29096
rect 19628 29084 19656 29112
rect 21266 29084 21272 29096
rect 19628 29056 21272 29084
rect 21266 29044 21272 29056
rect 21324 29044 21330 29096
rect 22830 29084 22836 29096
rect 22791 29056 22836 29084
rect 22830 29044 22836 29056
rect 22888 29044 22894 29096
rect 23017 29087 23075 29093
rect 23017 29053 23029 29087
rect 23063 29053 23075 29087
rect 23017 29047 23075 29053
rect 24029 29087 24087 29093
rect 24029 29053 24041 29087
rect 24075 29053 24087 29087
rect 24029 29047 24087 29053
rect 13814 29016 13820 29028
rect 12360 28988 12434 29016
rect 13727 28988 13820 29016
rect 8297 28951 8355 28957
rect 8297 28917 8309 28951
rect 8343 28948 8355 28951
rect 8386 28948 8392 28960
rect 8343 28920 8392 28948
rect 8343 28917 8355 28920
rect 8297 28911 8355 28917
rect 8386 28908 8392 28920
rect 8444 28948 8450 28960
rect 9582 28948 9588 28960
rect 8444 28920 9588 28948
rect 8444 28908 8450 28920
rect 9582 28908 9588 28920
rect 9640 28908 9646 28960
rect 12406 28948 12434 28988
rect 13740 28948 13768 28988
rect 13814 28976 13820 28988
rect 13872 29016 13878 29028
rect 14568 29016 14596 29044
rect 20073 29019 20131 29025
rect 20073 29016 20085 29019
rect 13872 28988 14596 29016
rect 19352 28988 20085 29016
rect 13872 28976 13878 28988
rect 14090 28948 14096 28960
rect 12406 28920 13768 28948
rect 14051 28920 14096 28948
rect 14090 28908 14096 28920
rect 14148 28908 14154 28960
rect 16298 28948 16304 28960
rect 16259 28920 16304 28948
rect 16298 28908 16304 28920
rect 16356 28908 16362 28960
rect 18711 28951 18769 28957
rect 18711 28917 18723 28951
rect 18757 28948 18769 28951
rect 19352 28948 19380 28988
rect 20073 28985 20085 28988
rect 20119 28985 20131 29019
rect 20073 28979 20131 28985
rect 22646 28976 22652 29028
rect 22704 29016 22710 29028
rect 23032 29016 23060 29047
rect 23566 29016 23572 29028
rect 22704 28988 23572 29016
rect 22704 28976 22710 28988
rect 23566 28976 23572 28988
rect 23624 28976 23630 29028
rect 24044 29016 24072 29047
rect 24118 29044 24124 29096
rect 24176 29084 24182 29096
rect 24854 29084 24860 29096
rect 24176 29056 24221 29084
rect 24815 29056 24860 29084
rect 24176 29044 24182 29056
rect 24854 29044 24860 29056
rect 24912 29044 24918 29096
rect 25130 29084 25136 29096
rect 25091 29056 25136 29084
rect 25130 29044 25136 29056
rect 25188 29044 25194 29096
rect 28442 29044 28448 29096
rect 28500 29084 28506 29096
rect 28626 29084 28632 29096
rect 28500 29056 28632 29084
rect 28500 29044 28506 29056
rect 28626 29044 28632 29056
rect 28684 29044 28690 29096
rect 28721 29087 28779 29093
rect 28721 29053 28733 29087
rect 28767 29053 28779 29087
rect 28721 29047 28779 29053
rect 26605 29019 26663 29025
rect 24044 28988 24900 29016
rect 18757 28920 19380 28948
rect 18757 28917 18769 28920
rect 18711 28911 18769 28917
rect 22094 28908 22100 28960
rect 22152 28948 22158 28960
rect 22373 28951 22431 28957
rect 22373 28948 22385 28951
rect 22152 28920 22385 28948
rect 22152 28908 22158 28920
rect 22373 28917 22385 28920
rect 22419 28917 22431 28951
rect 24872 28948 24900 28988
rect 26605 28985 26617 29019
rect 26651 29016 26663 29019
rect 26878 29016 26884 29028
rect 26651 28988 26884 29016
rect 26651 28985 26663 28988
rect 26605 28979 26663 28985
rect 26620 28948 26648 28979
rect 26878 28976 26884 28988
rect 26936 28976 26942 29028
rect 24872 28920 26648 28948
rect 28736 28948 28764 29047
rect 28810 29044 28816 29096
rect 28868 29084 28874 29096
rect 29012 29084 29040 29124
rect 29674 29121 29686 29124
rect 29720 29121 29732 29155
rect 29674 29115 29732 29121
rect 29822 29112 29828 29164
rect 29880 29152 29886 29164
rect 30208 29161 30236 29192
rect 31389 29189 31401 29223
rect 31435 29220 31447 29223
rect 32030 29220 32036 29232
rect 31435 29192 32036 29220
rect 31435 29189 31447 29192
rect 31389 29183 31447 29189
rect 32030 29180 32036 29192
rect 32088 29180 32094 29232
rect 34180 29223 34238 29229
rect 34180 29189 34192 29223
rect 34226 29220 34238 29223
rect 34900 29220 34928 29251
rect 34226 29192 34928 29220
rect 34226 29189 34238 29192
rect 34180 29183 34238 29189
rect 30101 29155 30159 29161
rect 30101 29152 30113 29155
rect 29880 29124 30113 29152
rect 29880 29112 29886 29124
rect 30101 29121 30113 29124
rect 30147 29121 30159 29155
rect 30101 29115 30159 29121
rect 30193 29155 30251 29161
rect 30193 29121 30205 29155
rect 30239 29121 30251 29155
rect 30193 29115 30251 29121
rect 31754 29112 31760 29164
rect 31812 29152 31818 29164
rect 32309 29155 32367 29161
rect 32309 29152 32321 29155
rect 31812 29124 32321 29152
rect 31812 29112 31818 29124
rect 32309 29121 32321 29124
rect 32355 29121 32367 29155
rect 32309 29115 32367 29121
rect 34514 29112 34520 29164
rect 34572 29152 34578 29164
rect 35069 29155 35127 29161
rect 35069 29152 35081 29155
rect 34572 29124 35081 29152
rect 34572 29112 34578 29124
rect 35069 29121 35081 29124
rect 35115 29121 35127 29155
rect 35069 29115 35127 29121
rect 28868 29056 29040 29084
rect 28868 29044 28874 29056
rect 30374 29044 30380 29096
rect 30432 29084 30438 29096
rect 31113 29087 31171 29093
rect 31113 29084 31125 29087
rect 30432 29056 31125 29084
rect 30432 29044 30438 29056
rect 31113 29053 31125 29056
rect 31159 29084 31171 29087
rect 33226 29084 33232 29096
rect 31159 29056 33232 29084
rect 31159 29053 31171 29056
rect 31113 29047 31171 29053
rect 33226 29044 33232 29056
rect 33284 29044 33290 29096
rect 34422 29084 34428 29096
rect 34383 29056 34428 29084
rect 34422 29044 34428 29056
rect 34480 29044 34486 29096
rect 29454 28948 29460 28960
rect 28736 28920 29460 28948
rect 22373 28911 22431 28917
rect 29454 28908 29460 28920
rect 29512 28908 29518 28960
rect 32490 28948 32496 28960
rect 32451 28920 32496 28948
rect 32490 28908 32496 28920
rect 32548 28908 32554 28960
rect 1104 28858 37628 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 37628 28858
rect 1104 28784 37628 28806
rect 10505 28747 10563 28753
rect 10505 28713 10517 28747
rect 10551 28744 10563 28747
rect 12618 28744 12624 28756
rect 10551 28716 12624 28744
rect 10551 28713 10563 28716
rect 10505 28707 10563 28713
rect 12618 28704 12624 28716
rect 12676 28704 12682 28756
rect 15562 28744 15568 28756
rect 15523 28716 15568 28744
rect 15562 28704 15568 28716
rect 15620 28704 15626 28756
rect 16114 28704 16120 28756
rect 16172 28744 16178 28756
rect 16853 28747 16911 28753
rect 16853 28744 16865 28747
rect 16172 28716 16865 28744
rect 16172 28704 16178 28716
rect 16853 28713 16865 28716
rect 16899 28713 16911 28747
rect 16853 28707 16911 28713
rect 25130 28704 25136 28756
rect 25188 28744 25194 28756
rect 25777 28747 25835 28753
rect 25777 28744 25789 28747
rect 25188 28716 25789 28744
rect 25188 28704 25194 28716
rect 25777 28713 25789 28716
rect 25823 28713 25835 28747
rect 26510 28744 26516 28756
rect 26471 28716 26516 28744
rect 25777 28707 25835 28713
rect 26510 28704 26516 28716
rect 26568 28704 26574 28756
rect 28994 28744 29000 28756
rect 28955 28716 29000 28744
rect 28994 28704 29000 28716
rect 29052 28704 29058 28756
rect 29086 28704 29092 28756
rect 29144 28744 29150 28756
rect 30285 28747 30343 28753
rect 30285 28744 30297 28747
rect 29144 28716 30297 28744
rect 29144 28704 29150 28716
rect 30285 28713 30297 28716
rect 30331 28713 30343 28747
rect 30285 28707 30343 28713
rect 31113 28747 31171 28753
rect 31113 28713 31125 28747
rect 31159 28744 31171 28747
rect 31294 28744 31300 28756
rect 31159 28716 31300 28744
rect 31159 28713 31171 28716
rect 31113 28707 31171 28713
rect 31294 28704 31300 28716
rect 31352 28704 31358 28756
rect 33873 28747 33931 28753
rect 33873 28713 33885 28747
rect 33919 28744 33931 28747
rect 34514 28744 34520 28756
rect 33919 28716 34520 28744
rect 33919 28713 33931 28716
rect 33873 28707 33931 28713
rect 34514 28704 34520 28716
rect 34572 28704 34578 28756
rect 9490 28636 9496 28688
rect 9548 28676 9554 28688
rect 14277 28679 14335 28685
rect 14277 28676 14289 28679
rect 9548 28648 9720 28676
rect 9548 28636 9554 28648
rect 8202 28568 8208 28620
rect 8260 28608 8266 28620
rect 8389 28611 8447 28617
rect 8389 28608 8401 28611
rect 8260 28580 8401 28608
rect 8260 28568 8266 28580
rect 8389 28577 8401 28580
rect 8435 28608 8447 28611
rect 9582 28608 9588 28620
rect 8435 28580 9444 28608
rect 9543 28580 9588 28608
rect 8435 28577 8447 28580
rect 8389 28571 8447 28577
rect 7193 28543 7251 28549
rect 7193 28509 7205 28543
rect 7239 28540 7251 28543
rect 7239 28512 7788 28540
rect 7239 28509 7251 28512
rect 7193 28503 7251 28509
rect 6822 28364 6828 28416
rect 6880 28404 6886 28416
rect 7760 28413 7788 28512
rect 8113 28475 8171 28481
rect 8113 28441 8125 28475
rect 8159 28472 8171 28475
rect 9416 28472 9444 28580
rect 9582 28568 9588 28580
rect 9640 28568 9646 28620
rect 9692 28617 9720 28648
rect 10336 28648 14289 28676
rect 9677 28611 9735 28617
rect 9677 28577 9689 28611
rect 9723 28577 9735 28611
rect 9677 28571 9735 28577
rect 10336 28549 10364 28648
rect 14277 28645 14289 28648
rect 14323 28645 14335 28679
rect 18138 28676 18144 28688
rect 14277 28639 14335 28645
rect 14936 28648 18144 28676
rect 11149 28611 11207 28617
rect 11149 28577 11161 28611
rect 11195 28577 11207 28611
rect 11149 28571 11207 28577
rect 10321 28543 10379 28549
rect 10321 28509 10333 28543
rect 10367 28509 10379 28543
rect 10321 28503 10379 28509
rect 11164 28472 11192 28571
rect 12526 28568 12532 28620
rect 12584 28608 12590 28620
rect 14936 28617 14964 28648
rect 18138 28636 18144 28648
rect 18196 28636 18202 28688
rect 25317 28679 25375 28685
rect 25317 28645 25329 28679
rect 25363 28645 25375 28679
rect 25317 28639 25375 28645
rect 12805 28611 12863 28617
rect 12805 28608 12817 28611
rect 12584 28580 12817 28608
rect 12584 28568 12590 28580
rect 12805 28577 12817 28580
rect 12851 28577 12863 28611
rect 14921 28611 14979 28617
rect 14921 28608 14933 28611
rect 12805 28571 12863 28577
rect 12912 28580 14933 28608
rect 12912 28540 12940 28580
rect 14921 28577 14933 28580
rect 14967 28577 14979 28611
rect 14921 28571 14979 28577
rect 17497 28611 17555 28617
rect 17497 28577 17509 28611
rect 17543 28608 17555 28611
rect 18230 28608 18236 28620
rect 17543 28580 18236 28608
rect 17543 28577 17555 28580
rect 17497 28571 17555 28577
rect 18230 28568 18236 28580
rect 18288 28568 18294 28620
rect 18414 28568 18420 28620
rect 18472 28608 18478 28620
rect 18601 28611 18659 28617
rect 18601 28608 18613 28611
rect 18472 28580 18613 28608
rect 18472 28568 18478 28580
rect 18601 28577 18613 28580
rect 18647 28577 18659 28611
rect 18601 28571 18659 28577
rect 18690 28568 18696 28620
rect 18748 28608 18754 28620
rect 18748 28580 18793 28608
rect 18748 28568 18754 28580
rect 18966 28568 18972 28620
rect 19024 28608 19030 28620
rect 20441 28611 20499 28617
rect 20441 28608 20453 28611
rect 19024 28580 20453 28608
rect 19024 28568 19030 28580
rect 20441 28577 20453 28580
rect 20487 28577 20499 28611
rect 20441 28571 20499 28577
rect 22189 28611 22247 28617
rect 22189 28577 22201 28611
rect 22235 28577 22247 28611
rect 22189 28571 22247 28577
rect 23845 28611 23903 28617
rect 23845 28577 23857 28611
rect 23891 28608 23903 28611
rect 24118 28608 24124 28620
rect 23891 28580 24124 28608
rect 23891 28577 23903 28580
rect 23845 28571 23903 28577
rect 12406 28512 12940 28540
rect 13725 28543 13783 28549
rect 12406 28472 12434 28512
rect 13725 28509 13737 28543
rect 13771 28540 13783 28543
rect 14182 28540 14188 28552
rect 13771 28512 14188 28540
rect 13771 28509 13783 28512
rect 13725 28503 13783 28509
rect 14182 28500 14188 28512
rect 14240 28500 14246 28552
rect 14642 28500 14648 28552
rect 14700 28500 14706 28552
rect 15470 28540 15476 28552
rect 15431 28512 15476 28540
rect 15470 28500 15476 28512
rect 15528 28500 15534 28552
rect 16301 28543 16359 28549
rect 16301 28509 16313 28543
rect 16347 28540 16359 28543
rect 16850 28540 16856 28552
rect 16347 28512 16856 28540
rect 16347 28509 16359 28512
rect 16301 28503 16359 28509
rect 16850 28500 16856 28512
rect 16908 28500 16914 28552
rect 17221 28543 17279 28549
rect 17221 28509 17233 28543
rect 17267 28540 17279 28543
rect 18432 28540 18460 28568
rect 17267 28512 18460 28540
rect 18708 28540 18736 28568
rect 19886 28540 19892 28552
rect 18708 28512 19892 28540
rect 17267 28509 17279 28512
rect 17221 28503 17279 28509
rect 19886 28500 19892 28512
rect 19944 28500 19950 28552
rect 19981 28543 20039 28549
rect 19981 28509 19993 28543
rect 20027 28509 20039 28543
rect 22204 28540 22232 28571
rect 24118 28568 24124 28580
rect 24176 28568 24182 28620
rect 24765 28611 24823 28617
rect 24765 28577 24777 28611
rect 24811 28608 24823 28611
rect 24946 28608 24952 28620
rect 24811 28580 24952 28608
rect 24811 28577 24823 28580
rect 24765 28571 24823 28577
rect 24946 28568 24952 28580
rect 25004 28608 25010 28620
rect 25130 28608 25136 28620
rect 25004 28580 25136 28608
rect 25004 28568 25010 28580
rect 25130 28568 25136 28580
rect 25188 28568 25194 28620
rect 22830 28540 22836 28552
rect 22204 28512 22836 28540
rect 19981 28503 20039 28509
rect 8159 28444 9168 28472
rect 9416 28444 12434 28472
rect 12529 28475 12587 28481
rect 8159 28441 8171 28444
rect 8113 28435 8171 28441
rect 7009 28407 7067 28413
rect 7009 28404 7021 28407
rect 6880 28376 7021 28404
rect 6880 28364 6886 28376
rect 7009 28373 7021 28376
rect 7055 28373 7067 28407
rect 7009 28367 7067 28373
rect 7745 28407 7803 28413
rect 7745 28373 7757 28407
rect 7791 28373 7803 28407
rect 7745 28367 7803 28373
rect 8205 28407 8263 28413
rect 8205 28373 8217 28407
rect 8251 28404 8263 28407
rect 8294 28404 8300 28416
rect 8251 28376 8300 28404
rect 8251 28373 8263 28376
rect 8205 28367 8263 28373
rect 8294 28364 8300 28376
rect 8352 28364 8358 28416
rect 9140 28413 9168 28444
rect 12529 28441 12541 28475
rect 12575 28472 12587 28475
rect 14660 28472 14688 28500
rect 14826 28472 14832 28484
rect 12575 28444 14832 28472
rect 12575 28441 12587 28444
rect 12529 28435 12587 28441
rect 14826 28432 14832 28444
rect 14884 28432 14890 28484
rect 19996 28472 20024 28503
rect 22830 28500 22836 28512
rect 22888 28540 22894 28552
rect 23569 28543 23627 28549
rect 23569 28540 23581 28543
rect 22888 28512 23581 28540
rect 22888 28500 22894 28512
rect 23569 28509 23581 28512
rect 23615 28540 23627 28543
rect 24857 28543 24915 28549
rect 24857 28540 24869 28543
rect 23615 28512 24869 28540
rect 23615 28509 23627 28512
rect 23569 28503 23627 28509
rect 24857 28509 24869 28512
rect 24903 28509 24915 28543
rect 25332 28540 25360 28639
rect 26878 28636 26884 28688
rect 26936 28676 26942 28688
rect 26936 28648 28856 28676
rect 26936 28636 26942 28648
rect 28350 28568 28356 28620
rect 28408 28608 28414 28620
rect 28537 28611 28595 28617
rect 28537 28608 28549 28611
rect 28408 28580 28549 28608
rect 28408 28568 28414 28580
rect 28537 28577 28549 28580
rect 28583 28577 28595 28611
rect 28537 28571 28595 28577
rect 28629 28611 28687 28617
rect 28629 28577 28641 28611
rect 28675 28608 28687 28611
rect 28718 28608 28724 28620
rect 28675 28580 28724 28608
rect 28675 28577 28687 28580
rect 28629 28571 28687 28577
rect 28718 28568 28724 28580
rect 28776 28568 28782 28620
rect 28828 28608 28856 28648
rect 29178 28636 29184 28688
rect 29236 28676 29242 28688
rect 29236 28648 30052 28676
rect 29236 28636 29242 28648
rect 29638 28608 29644 28620
rect 28828 28580 29644 28608
rect 25961 28543 26019 28549
rect 25961 28540 25973 28543
rect 25332 28512 25973 28540
rect 24857 28503 24915 28509
rect 25961 28509 25973 28512
rect 26007 28509 26019 28543
rect 26602 28540 26608 28552
rect 26563 28512 26608 28540
rect 25961 28503 26019 28509
rect 26602 28500 26608 28512
rect 26660 28500 26666 28552
rect 28258 28540 28264 28552
rect 28219 28512 28264 28540
rect 28258 28500 28264 28512
rect 28316 28500 28322 28552
rect 28828 28549 28856 28580
rect 29638 28568 29644 28580
rect 29696 28568 29702 28620
rect 28445 28543 28503 28549
rect 28445 28509 28457 28543
rect 28491 28509 28503 28543
rect 28445 28503 28503 28509
rect 28813 28543 28871 28549
rect 28813 28509 28825 28543
rect 28859 28509 28871 28543
rect 28813 28503 28871 28509
rect 20717 28475 20775 28481
rect 19996 28444 20576 28472
rect 20548 28416 20576 28444
rect 20717 28441 20729 28475
rect 20763 28472 20775 28475
rect 20806 28472 20812 28484
rect 20763 28444 20812 28472
rect 20763 28441 20775 28444
rect 20717 28435 20775 28441
rect 20806 28432 20812 28444
rect 20864 28432 20870 28484
rect 23474 28472 23480 28484
rect 21942 28444 23480 28472
rect 23474 28432 23480 28444
rect 23532 28432 23538 28484
rect 24949 28475 25007 28481
rect 24949 28441 24961 28475
rect 24995 28472 25007 28475
rect 26878 28472 26884 28484
rect 24995 28444 26884 28472
rect 24995 28441 25007 28444
rect 24949 28435 25007 28441
rect 26878 28432 26884 28444
rect 26936 28432 26942 28484
rect 28460 28472 28488 28503
rect 28902 28500 28908 28552
rect 28960 28540 28966 28552
rect 29733 28543 29791 28549
rect 29733 28540 29745 28543
rect 28960 28512 29745 28540
rect 28960 28500 28966 28512
rect 29733 28509 29745 28512
rect 29779 28509 29791 28543
rect 29733 28503 29791 28509
rect 29822 28500 29828 28552
rect 29880 28540 29886 28552
rect 30024 28549 30052 28648
rect 33226 28608 33232 28620
rect 33187 28580 33232 28608
rect 33226 28568 33232 28580
rect 33284 28568 33290 28620
rect 30009 28543 30067 28549
rect 29880 28512 29925 28540
rect 29880 28500 29886 28512
rect 30009 28509 30021 28543
rect 30055 28509 30067 28543
rect 30009 28503 30067 28509
rect 30101 28543 30159 28549
rect 30101 28509 30113 28543
rect 30147 28509 30159 28543
rect 30101 28503 30159 28509
rect 28534 28472 28540 28484
rect 28447 28444 28540 28472
rect 28534 28432 28540 28444
rect 28592 28472 28598 28484
rect 29270 28472 29276 28484
rect 28592 28444 29276 28472
rect 28592 28432 28598 28444
rect 29270 28432 29276 28444
rect 29328 28432 29334 28484
rect 29454 28432 29460 28484
rect 29512 28472 29518 28484
rect 30116 28472 30144 28503
rect 31938 28500 31944 28552
rect 31996 28540 32002 28552
rect 32493 28543 32551 28549
rect 32493 28540 32505 28543
rect 31996 28512 32505 28540
rect 31996 28500 32002 28512
rect 32493 28509 32505 28512
rect 32539 28509 32551 28543
rect 32493 28503 32551 28509
rect 33134 28500 33140 28552
rect 33192 28540 33198 28552
rect 33413 28543 33471 28549
rect 33413 28540 33425 28543
rect 33192 28512 33425 28540
rect 33192 28500 33198 28512
rect 33413 28509 33425 28512
rect 33459 28509 33471 28543
rect 33413 28503 33471 28509
rect 34885 28543 34943 28549
rect 34885 28509 34897 28543
rect 34931 28509 34943 28543
rect 35066 28540 35072 28552
rect 35027 28512 35072 28540
rect 34885 28503 34943 28509
rect 29512 28444 30144 28472
rect 32248 28475 32306 28481
rect 29512 28432 29518 28444
rect 32248 28441 32260 28475
rect 32294 28472 32306 28475
rect 32398 28472 32404 28484
rect 32294 28444 32404 28472
rect 32294 28441 32306 28444
rect 32248 28435 32306 28441
rect 32398 28432 32404 28444
rect 32456 28432 32462 28484
rect 34900 28472 34928 28503
rect 35066 28500 35072 28512
rect 35124 28500 35130 28552
rect 35434 28500 35440 28552
rect 35492 28540 35498 28552
rect 35713 28543 35771 28549
rect 35713 28540 35725 28543
rect 35492 28512 35725 28540
rect 35492 28500 35498 28512
rect 35713 28509 35725 28512
rect 35759 28509 35771 28543
rect 35713 28503 35771 28509
rect 32508 28444 34928 28472
rect 9125 28407 9183 28413
rect 9125 28373 9137 28407
rect 9171 28373 9183 28407
rect 9125 28367 9183 28373
rect 9214 28364 9220 28416
rect 9272 28404 9278 28416
rect 9493 28407 9551 28413
rect 9493 28404 9505 28407
rect 9272 28376 9505 28404
rect 9272 28364 9278 28376
rect 9493 28373 9505 28376
rect 9539 28373 9551 28407
rect 11238 28404 11244 28416
rect 11199 28376 11244 28404
rect 9493 28367 9551 28373
rect 11238 28364 11244 28376
rect 11296 28364 11302 28416
rect 11330 28364 11336 28416
rect 11388 28404 11394 28416
rect 11701 28407 11759 28413
rect 11388 28376 11433 28404
rect 11388 28364 11394 28376
rect 11701 28373 11713 28407
rect 11747 28404 11759 28407
rect 11882 28404 11888 28416
rect 11747 28376 11888 28404
rect 11747 28373 11759 28376
rect 11701 28367 11759 28373
rect 11882 28364 11888 28376
rect 11940 28364 11946 28416
rect 13538 28404 13544 28416
rect 13499 28376 13544 28404
rect 13538 28364 13544 28376
rect 13596 28364 13602 28416
rect 14642 28404 14648 28416
rect 14603 28376 14648 28404
rect 14642 28364 14648 28376
rect 14700 28364 14706 28416
rect 14734 28364 14740 28416
rect 14792 28404 14798 28416
rect 16114 28404 16120 28416
rect 14792 28376 14837 28404
rect 16075 28376 16120 28404
rect 14792 28364 14798 28376
rect 16114 28364 16120 28376
rect 16172 28364 16178 28416
rect 17313 28407 17371 28413
rect 17313 28373 17325 28407
rect 17359 28404 17371 28407
rect 17586 28404 17592 28416
rect 17359 28376 17592 28404
rect 17359 28373 17371 28376
rect 17313 28367 17371 28373
rect 17586 28364 17592 28376
rect 17644 28364 17650 28416
rect 18046 28364 18052 28416
rect 18104 28404 18110 28416
rect 18141 28407 18199 28413
rect 18141 28404 18153 28407
rect 18104 28376 18153 28404
rect 18104 28364 18110 28376
rect 18141 28373 18153 28376
rect 18187 28373 18199 28407
rect 18141 28367 18199 28373
rect 18414 28364 18420 28416
rect 18472 28404 18478 28416
rect 18509 28407 18567 28413
rect 18509 28404 18521 28407
rect 18472 28376 18521 28404
rect 18472 28364 18478 28376
rect 18509 28373 18521 28376
rect 18555 28373 18567 28407
rect 18509 28367 18567 28373
rect 19889 28407 19947 28413
rect 19889 28373 19901 28407
rect 19935 28404 19947 28407
rect 19978 28404 19984 28416
rect 19935 28376 19984 28404
rect 19935 28373 19947 28376
rect 19889 28367 19947 28373
rect 19978 28364 19984 28376
rect 20036 28364 20042 28416
rect 20530 28364 20536 28416
rect 20588 28364 20594 28416
rect 23198 28404 23204 28416
rect 23159 28376 23204 28404
rect 23198 28364 23204 28376
rect 23256 28364 23262 28416
rect 23661 28407 23719 28413
rect 23661 28373 23673 28407
rect 23707 28404 23719 28407
rect 24578 28404 24584 28416
rect 23707 28376 24584 28404
rect 23707 28373 23719 28376
rect 23661 28367 23719 28373
rect 24578 28364 24584 28376
rect 24636 28364 24642 28416
rect 29914 28364 29920 28416
rect 29972 28404 29978 28416
rect 31018 28404 31024 28416
rect 29972 28376 31024 28404
rect 29972 28364 29978 28376
rect 31018 28364 31024 28376
rect 31076 28364 31082 28416
rect 31202 28364 31208 28416
rect 31260 28404 31266 28416
rect 32508 28404 32536 28444
rect 31260 28376 32536 28404
rect 31260 28364 31266 28376
rect 33410 28364 33416 28416
rect 33468 28404 33474 28416
rect 33505 28407 33563 28413
rect 33505 28404 33517 28407
rect 33468 28376 33517 28404
rect 33468 28364 33474 28376
rect 33505 28373 33517 28376
rect 33551 28373 33563 28407
rect 33505 28367 33563 28373
rect 34606 28364 34612 28416
rect 34664 28404 34670 28416
rect 34977 28407 35035 28413
rect 34977 28404 34989 28407
rect 34664 28376 34989 28404
rect 34664 28364 34670 28376
rect 34977 28373 34989 28376
rect 35023 28373 35035 28407
rect 34977 28367 35035 28373
rect 35158 28364 35164 28416
rect 35216 28404 35222 28416
rect 35529 28407 35587 28413
rect 35529 28404 35541 28407
rect 35216 28376 35541 28404
rect 35216 28364 35222 28376
rect 35529 28373 35541 28376
rect 35575 28373 35587 28407
rect 35529 28367 35587 28373
rect 1104 28314 37628 28336
rect 1104 28262 4874 28314
rect 4926 28262 4938 28314
rect 4990 28262 5002 28314
rect 5054 28262 5066 28314
rect 5118 28262 5130 28314
rect 5182 28262 35594 28314
rect 35646 28262 35658 28314
rect 35710 28262 35722 28314
rect 35774 28262 35786 28314
rect 35838 28262 35850 28314
rect 35902 28262 37628 28314
rect 1104 28240 37628 28262
rect 7098 28200 7104 28212
rect 6564 28172 7104 28200
rect 1765 28067 1823 28073
rect 1765 28033 1777 28067
rect 1811 28064 1823 28067
rect 1854 28064 1860 28076
rect 1811 28036 1860 28064
rect 1811 28033 1823 28036
rect 1765 28027 1823 28033
rect 1854 28024 1860 28036
rect 1912 28024 1918 28076
rect 6564 28073 6592 28172
rect 7098 28160 7104 28172
rect 7156 28200 7162 28212
rect 8294 28200 8300 28212
rect 7156 28172 8156 28200
rect 8255 28172 8300 28200
rect 7156 28160 7162 28172
rect 6822 28132 6828 28144
rect 6783 28104 6828 28132
rect 6822 28092 6828 28104
rect 6880 28092 6886 28144
rect 7282 28092 7288 28144
rect 7340 28092 7346 28144
rect 6549 28067 6607 28073
rect 6549 28033 6561 28067
rect 6595 28033 6607 28067
rect 6549 28027 6607 28033
rect 8128 27996 8156 28172
rect 8294 28160 8300 28172
rect 8352 28160 8358 28212
rect 11149 28203 11207 28209
rect 11149 28169 11161 28203
rect 11195 28200 11207 28203
rect 11238 28200 11244 28212
rect 11195 28172 11244 28200
rect 11195 28169 11207 28172
rect 11149 28163 11207 28169
rect 11238 28160 11244 28172
rect 11296 28160 11302 28212
rect 11330 28160 11336 28212
rect 11388 28200 11394 28212
rect 12345 28203 12403 28209
rect 12345 28200 12357 28203
rect 11388 28172 12357 28200
rect 11388 28160 11394 28172
rect 12345 28169 12357 28172
rect 12391 28169 12403 28203
rect 14182 28200 14188 28212
rect 14143 28172 14188 28200
rect 12345 28163 12403 28169
rect 14182 28160 14188 28172
rect 14240 28160 14246 28212
rect 14642 28160 14648 28212
rect 14700 28200 14706 28212
rect 15381 28203 15439 28209
rect 15381 28200 15393 28203
rect 14700 28172 15393 28200
rect 14700 28160 14706 28172
rect 15381 28169 15393 28172
rect 15427 28169 15439 28203
rect 16850 28200 16856 28212
rect 16811 28172 16856 28200
rect 15381 28163 15439 28169
rect 16850 28160 16856 28172
rect 16908 28160 16914 28212
rect 18233 28203 18291 28209
rect 18233 28169 18245 28203
rect 18279 28200 18291 28203
rect 18279 28172 19012 28200
rect 18279 28169 18291 28172
rect 18233 28163 18291 28169
rect 8849 28135 8907 28141
rect 8849 28101 8861 28135
rect 8895 28132 8907 28135
rect 12713 28135 12771 28141
rect 8895 28104 10166 28132
rect 8895 28101 8907 28104
rect 8849 28095 8907 28101
rect 12713 28101 12725 28135
rect 12759 28132 12771 28135
rect 14090 28132 14096 28144
rect 12759 28104 14096 28132
rect 12759 28101 12771 28104
rect 12713 28095 12771 28101
rect 14090 28092 14096 28104
rect 14148 28132 14154 28144
rect 14734 28132 14740 28144
rect 14148 28104 14740 28132
rect 14148 28092 14154 28104
rect 8754 28064 8760 28076
rect 8715 28036 8760 28064
rect 8754 28024 8760 28036
rect 8812 28024 8818 28076
rect 9401 28067 9459 28073
rect 9401 28033 9413 28067
rect 9447 28033 9459 28067
rect 11882 28064 11888 28076
rect 11843 28036 11888 28064
rect 9401 28027 9459 28033
rect 9306 27996 9312 28008
rect 8128 27968 9312 27996
rect 9306 27956 9312 27968
rect 9364 27996 9370 28008
rect 9416 27996 9444 28027
rect 11882 28024 11888 28036
rect 11940 28024 11946 28076
rect 12805 28067 12863 28073
rect 12805 28033 12817 28067
rect 12851 28064 12863 28067
rect 13078 28064 13084 28076
rect 12851 28036 13084 28064
rect 12851 28033 12863 28036
rect 12805 28027 12863 28033
rect 13078 28024 13084 28036
rect 13136 28024 13142 28076
rect 13541 28067 13599 28073
rect 13541 28033 13553 28067
rect 13587 28064 13599 28067
rect 13722 28064 13728 28076
rect 13587 28036 13728 28064
rect 13587 28033 13599 28036
rect 13541 28027 13599 28033
rect 13722 28024 13728 28036
rect 13780 28024 13786 28076
rect 14660 28073 14688 28104
rect 14734 28092 14740 28104
rect 14792 28092 14798 28144
rect 15749 28135 15807 28141
rect 15749 28101 15761 28135
rect 15795 28132 15807 28135
rect 16298 28132 16304 28144
rect 15795 28104 16304 28132
rect 15795 28101 15807 28104
rect 15749 28095 15807 28101
rect 16298 28092 16304 28104
rect 16356 28132 16362 28144
rect 17313 28135 17371 28141
rect 17313 28132 17325 28135
rect 16356 28104 17325 28132
rect 16356 28092 16362 28104
rect 17313 28101 17325 28104
rect 17359 28101 17371 28135
rect 18690 28132 18696 28144
rect 17313 28095 17371 28101
rect 18616 28104 18696 28132
rect 14553 28067 14611 28073
rect 14553 28033 14565 28067
rect 14599 28033 14611 28067
rect 14553 28027 14611 28033
rect 14645 28067 14703 28073
rect 14645 28033 14657 28067
rect 14691 28033 14703 28067
rect 17221 28067 17279 28073
rect 14645 28027 14703 28033
rect 14844 28036 17172 28064
rect 9364 27968 9444 27996
rect 9677 27999 9735 28005
rect 9364 27956 9370 27968
rect 9677 27965 9689 27999
rect 9723 27996 9735 27999
rect 9723 27968 11744 27996
rect 9723 27965 9735 27968
rect 9677 27959 9735 27965
rect 11716 27937 11744 27968
rect 12710 27956 12716 28008
rect 12768 27996 12774 28008
rect 12897 27999 12955 28005
rect 12897 27996 12909 27999
rect 12768 27968 12909 27996
rect 12768 27956 12774 27968
rect 12897 27965 12909 27968
rect 12943 27965 12955 27999
rect 12897 27959 12955 27965
rect 11701 27931 11759 27937
rect 11701 27897 11713 27931
rect 11747 27897 11759 27931
rect 14568 27928 14596 28027
rect 14844 28005 14872 28036
rect 14829 27999 14887 28005
rect 14829 27965 14841 27999
rect 14875 27965 14887 27999
rect 14829 27959 14887 27965
rect 15841 27999 15899 28005
rect 15841 27965 15853 27999
rect 15887 27965 15899 27999
rect 15841 27959 15899 27965
rect 16025 27999 16083 28005
rect 16025 27965 16037 27999
rect 16071 27965 16083 27999
rect 17144 27996 17172 28036
rect 17221 28033 17233 28067
rect 17267 28064 17279 28067
rect 17586 28064 17592 28076
rect 17267 28036 17592 28064
rect 17267 28033 17279 28036
rect 17221 28027 17279 28033
rect 17586 28024 17592 28036
rect 17644 28024 17650 28076
rect 18046 28064 18052 28076
rect 18007 28036 18052 28064
rect 18046 28024 18052 28036
rect 18104 28024 18110 28076
rect 17405 27999 17463 28005
rect 17405 27996 17417 27999
rect 17144 27968 17417 27996
rect 16025 27959 16083 27965
rect 17405 27965 17417 27968
rect 17451 27996 17463 27999
rect 18616 27996 18644 28104
rect 18690 28092 18696 28104
rect 18748 28092 18754 28144
rect 18984 28141 19012 28172
rect 20806 28160 20812 28212
rect 20864 28200 20870 28212
rect 20901 28203 20959 28209
rect 20901 28200 20913 28203
rect 20864 28172 20913 28200
rect 20864 28160 20870 28172
rect 20901 28169 20913 28172
rect 20947 28169 20959 28203
rect 20901 28163 20959 28169
rect 28258 28160 28264 28212
rect 28316 28200 28322 28212
rect 28721 28203 28779 28209
rect 28721 28200 28733 28203
rect 28316 28172 28733 28200
rect 28316 28160 28322 28172
rect 28721 28169 28733 28172
rect 28767 28169 28779 28203
rect 28721 28163 28779 28169
rect 29825 28203 29883 28209
rect 29825 28169 29837 28203
rect 29871 28200 29883 28203
rect 29914 28200 29920 28212
rect 29871 28172 29920 28200
rect 29871 28169 29883 28172
rect 29825 28163 29883 28169
rect 29914 28160 29920 28172
rect 29972 28160 29978 28212
rect 30742 28200 30748 28212
rect 30024 28172 30748 28200
rect 18969 28135 19027 28141
rect 18969 28101 18981 28135
rect 19015 28101 19027 28135
rect 18969 28095 19027 28101
rect 19978 28092 19984 28144
rect 20036 28092 20042 28144
rect 22278 28092 22284 28144
rect 22336 28132 22342 28144
rect 22336 28104 23060 28132
rect 22336 28092 22342 28104
rect 23032 28076 23060 28104
rect 24762 28092 24768 28144
rect 24820 28132 24826 28144
rect 25317 28135 25375 28141
rect 25317 28132 25329 28135
rect 24820 28104 25329 28132
rect 24820 28092 24826 28104
rect 25317 28101 25329 28104
rect 25363 28101 25375 28135
rect 25317 28095 25375 28101
rect 21085 28067 21143 28073
rect 21085 28033 21097 28067
rect 21131 28064 21143 28067
rect 22094 28064 22100 28076
rect 21131 28036 22100 28064
rect 21131 28033 21143 28036
rect 21085 28027 21143 28033
rect 22094 28024 22100 28036
rect 22152 28024 22158 28076
rect 22186 28024 22192 28076
rect 22244 28064 22250 28076
rect 23014 28064 23020 28076
rect 22244 28036 22289 28064
rect 22975 28036 23020 28064
rect 22244 28024 22250 28036
rect 23014 28024 23020 28036
rect 23072 28024 23078 28076
rect 24210 28064 24216 28076
rect 24171 28036 24216 28064
rect 24210 28024 24216 28036
rect 24268 28024 24274 28076
rect 24305 28067 24363 28073
rect 24305 28033 24317 28067
rect 24351 28064 24363 28067
rect 25409 28067 25467 28073
rect 25409 28064 25421 28067
rect 24351 28036 25421 28064
rect 24351 28033 24363 28036
rect 24305 28027 24363 28033
rect 25409 28033 25421 28036
rect 25455 28033 25467 28067
rect 25409 28027 25467 28033
rect 26421 28067 26479 28073
rect 26421 28033 26433 28067
rect 26467 28064 26479 28067
rect 26602 28064 26608 28076
rect 26467 28036 26608 28064
rect 26467 28033 26479 28036
rect 26421 28027 26479 28033
rect 17451 27968 18644 27996
rect 18693 27999 18751 28005
rect 17451 27965 17463 27968
rect 17405 27959 17463 27965
rect 18693 27965 18705 27999
rect 18739 27996 18751 27999
rect 23293 27999 23351 28005
rect 18739 27968 18828 27996
rect 18739 27965 18751 27968
rect 18693 27959 18751 27965
rect 15010 27928 15016 27940
rect 14568 27900 15016 27928
rect 11701 27891 11759 27897
rect 15010 27888 15016 27900
rect 15068 27928 15074 27940
rect 15856 27928 15884 27959
rect 15068 27900 15884 27928
rect 16040 27928 16068 27959
rect 18230 27928 18236 27940
rect 16040 27900 18236 27928
rect 15068 27888 15074 27900
rect 18230 27888 18236 27900
rect 18288 27888 18294 27940
rect 1578 27860 1584 27872
rect 1539 27832 1584 27860
rect 1578 27820 1584 27832
rect 1636 27820 1642 27872
rect 13630 27860 13636 27872
rect 13591 27832 13636 27860
rect 13630 27820 13636 27832
rect 13688 27820 13694 27872
rect 18800 27860 18828 27968
rect 23293 27965 23305 27999
rect 23339 27996 23351 27999
rect 24118 27996 24124 28008
rect 23339 27968 24124 27996
rect 23339 27965 23351 27968
rect 23293 27959 23351 27965
rect 24118 27956 24124 27968
rect 24176 27996 24182 28008
rect 24397 27999 24455 28005
rect 24397 27996 24409 27999
rect 24176 27968 24409 27996
rect 24176 27956 24182 27968
rect 24397 27965 24409 27968
rect 24443 27965 24455 27999
rect 25130 27996 25136 28008
rect 25091 27968 25136 27996
rect 24397 27959 24455 27965
rect 25130 27956 25136 27968
rect 25188 27956 25194 28008
rect 25424 27996 25452 28027
rect 26602 28024 26608 28036
rect 26660 28024 26666 28076
rect 27893 28067 27951 28073
rect 27893 28033 27905 28067
rect 27939 28064 27951 28067
rect 28810 28064 28816 28076
rect 27939 28036 28816 28064
rect 27939 28033 27951 28036
rect 27893 28027 27951 28033
rect 27908 27996 27936 28027
rect 28810 28024 28816 28036
rect 28868 28064 28874 28076
rect 30024 28073 30052 28172
rect 30742 28160 30748 28172
rect 30800 28200 30806 28212
rect 33502 28200 33508 28212
rect 30800 28172 33508 28200
rect 30800 28160 30806 28172
rect 33502 28160 33508 28172
rect 33560 28200 33566 28212
rect 34057 28203 34115 28209
rect 33560 28172 34008 28200
rect 33560 28160 33566 28172
rect 32401 28135 32459 28141
rect 32401 28101 32413 28135
rect 32447 28132 32459 28135
rect 32490 28132 32496 28144
rect 32447 28104 32496 28132
rect 32447 28101 32459 28104
rect 32401 28095 32459 28101
rect 32490 28092 32496 28104
rect 32548 28092 32554 28144
rect 32950 28092 32956 28144
rect 33008 28132 33014 28144
rect 33008 28104 33548 28132
rect 33008 28092 33014 28104
rect 28997 28067 29055 28073
rect 28997 28064 29009 28067
rect 28868 28036 29009 28064
rect 28868 28024 28874 28036
rect 28997 28033 29009 28036
rect 29043 28033 29055 28067
rect 28997 28027 29055 28033
rect 29273 28067 29331 28073
rect 29273 28033 29285 28067
rect 29319 28033 29331 28067
rect 29273 28027 29331 28033
rect 29733 28067 29791 28073
rect 29733 28033 29745 28067
rect 29779 28033 29791 28067
rect 29733 28027 29791 28033
rect 30009 28067 30067 28073
rect 30009 28033 30021 28067
rect 30055 28033 30067 28067
rect 30009 28027 30067 28033
rect 30193 28067 30251 28073
rect 30193 28033 30205 28067
rect 30239 28064 30251 28067
rect 30653 28067 30711 28073
rect 30653 28064 30665 28067
rect 30239 28036 30665 28064
rect 30239 28033 30251 28036
rect 30193 28027 30251 28033
rect 30653 28033 30665 28036
rect 30699 28033 30711 28067
rect 30653 28027 30711 28033
rect 31021 28067 31079 28073
rect 31021 28033 31033 28067
rect 31067 28064 31079 28067
rect 31110 28064 31116 28076
rect 31067 28036 31116 28064
rect 31067 28033 31079 28036
rect 31021 28027 31079 28033
rect 25424 27968 27936 27996
rect 27985 27999 28043 28005
rect 27985 27965 27997 27999
rect 28031 27965 28043 27999
rect 27985 27959 28043 27965
rect 28261 27999 28319 28005
rect 28261 27965 28273 27999
rect 28307 27996 28319 27999
rect 28902 27996 28908 28008
rect 28307 27968 28908 27996
rect 28307 27965 28319 27968
rect 28261 27959 28319 27965
rect 28000 27928 28028 27959
rect 28902 27956 28908 27968
rect 28960 27956 28966 28008
rect 29288 27928 29316 28027
rect 29748 27996 29776 28027
rect 31110 28024 31116 28036
rect 31168 28024 31174 28076
rect 31205 28067 31263 28073
rect 31205 28033 31217 28067
rect 31251 28064 31263 28067
rect 31570 28064 31576 28076
rect 31251 28036 31576 28064
rect 31251 28033 31263 28036
rect 31205 28027 31263 28033
rect 31570 28024 31576 28036
rect 31628 28064 31634 28076
rect 33520 28073 33548 28104
rect 33980 28073 34008 28172
rect 34057 28169 34069 28203
rect 34103 28200 34115 28203
rect 35066 28200 35072 28212
rect 34103 28172 35072 28200
rect 34103 28169 34115 28172
rect 34057 28163 34115 28169
rect 35066 28160 35072 28172
rect 35124 28160 35130 28212
rect 34422 28132 34428 28144
rect 34072 28104 34428 28132
rect 33413 28067 33471 28073
rect 33413 28064 33425 28067
rect 31628 28036 33425 28064
rect 31628 28024 31634 28036
rect 33413 28033 33425 28036
rect 33459 28033 33471 28067
rect 33413 28027 33471 28033
rect 33505 28067 33563 28073
rect 33505 28033 33517 28067
rect 33551 28033 33563 28067
rect 33505 28027 33563 28033
rect 33965 28067 34023 28073
rect 33965 28033 33977 28067
rect 34011 28033 34023 28067
rect 33965 28027 34023 28033
rect 30558 27996 30564 28008
rect 29748 27968 30564 27996
rect 30558 27956 30564 27968
rect 30616 27996 30622 28008
rect 31386 27996 31392 28008
rect 30616 27968 31392 27996
rect 30616 27956 30622 27968
rect 31386 27956 31392 27968
rect 31444 27956 31450 28008
rect 31938 27956 31944 28008
rect 31996 27996 32002 28008
rect 34072 27996 34100 28104
rect 34422 28092 34428 28104
rect 34480 28132 34486 28144
rect 35158 28132 35164 28144
rect 34480 28104 34928 28132
rect 35119 28104 35164 28132
rect 34480 28092 34486 28104
rect 34149 28067 34207 28073
rect 34149 28033 34161 28067
rect 34195 28033 34207 28067
rect 34149 28027 34207 28033
rect 31996 27968 34100 27996
rect 31996 27956 32002 27968
rect 30466 27928 30472 27940
rect 28000 27900 30472 27928
rect 30466 27888 30472 27900
rect 30524 27888 30530 27940
rect 31021 27931 31079 27937
rect 31021 27897 31033 27931
rect 31067 27928 31079 27931
rect 33318 27928 33324 27940
rect 31067 27900 33324 27928
rect 31067 27897 31079 27900
rect 31021 27891 31079 27897
rect 33318 27888 33324 27900
rect 33376 27888 33382 27940
rect 18966 27860 18972 27872
rect 18800 27832 18972 27860
rect 18966 27820 18972 27832
rect 19024 27860 19030 27872
rect 19702 27860 19708 27872
rect 19024 27832 19708 27860
rect 19024 27820 19030 27832
rect 19702 27820 19708 27832
rect 19760 27820 19766 27872
rect 20438 27860 20444 27872
rect 20399 27832 20444 27860
rect 20438 27820 20444 27832
rect 20496 27820 20502 27872
rect 22094 27820 22100 27872
rect 22152 27860 22158 27872
rect 23842 27860 23848 27872
rect 22152 27832 22197 27860
rect 23803 27832 23848 27860
rect 22152 27820 22158 27832
rect 23842 27820 23848 27832
rect 23900 27820 23906 27872
rect 25777 27863 25835 27869
rect 25777 27829 25789 27863
rect 25823 27860 25835 27863
rect 26142 27860 26148 27872
rect 25823 27832 26148 27860
rect 25823 27829 25835 27832
rect 25777 27823 25835 27829
rect 26142 27820 26148 27832
rect 26200 27820 26206 27872
rect 26513 27863 26571 27869
rect 26513 27829 26525 27863
rect 26559 27860 26571 27863
rect 27522 27860 27528 27872
rect 26559 27832 27528 27860
rect 26559 27829 26571 27832
rect 26513 27823 26571 27829
rect 27522 27820 27528 27832
rect 27580 27820 27586 27872
rect 29178 27860 29184 27872
rect 29091 27832 29184 27860
rect 29178 27820 29184 27832
rect 29236 27860 29242 27872
rect 29822 27860 29828 27872
rect 29236 27832 29828 27860
rect 29236 27820 29242 27832
rect 29822 27820 29828 27832
rect 29880 27820 29886 27872
rect 32030 27820 32036 27872
rect 32088 27860 32094 27872
rect 32493 27863 32551 27869
rect 32493 27860 32505 27863
rect 32088 27832 32505 27860
rect 32088 27820 32094 27832
rect 32493 27829 32505 27832
rect 32539 27860 32551 27863
rect 34164 27860 34192 28027
rect 34900 28005 34928 28104
rect 35158 28092 35164 28104
rect 35216 28092 35222 28144
rect 36170 28092 36176 28144
rect 36228 28092 36234 28144
rect 34885 27999 34943 28005
rect 34885 27965 34897 27999
rect 34931 27965 34943 27999
rect 34885 27959 34943 27965
rect 36630 27860 36636 27872
rect 32539 27832 34192 27860
rect 36591 27832 36636 27860
rect 32539 27829 32551 27832
rect 32493 27823 32551 27829
rect 36630 27820 36636 27832
rect 36688 27820 36694 27872
rect 1104 27770 37628 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 37628 27770
rect 1104 27696 37628 27718
rect 16114 27665 16120 27668
rect 16104 27659 16120 27665
rect 16104 27625 16116 27659
rect 16104 27619 16120 27625
rect 16114 27616 16120 27619
rect 16172 27616 16178 27668
rect 22186 27616 22192 27668
rect 22244 27656 22250 27668
rect 22244 27628 23612 27656
rect 22244 27616 22250 27628
rect 7282 27588 7288 27600
rect 7243 27560 7288 27588
rect 7282 27548 7288 27560
rect 7340 27548 7346 27600
rect 14550 27548 14556 27600
rect 14608 27588 14614 27600
rect 14608 27560 15884 27588
rect 14608 27548 14614 27560
rect 8202 27480 8208 27532
rect 8260 27520 8266 27532
rect 8389 27523 8447 27529
rect 8389 27520 8401 27523
rect 8260 27492 8401 27520
rect 8260 27480 8266 27492
rect 8389 27489 8401 27492
rect 8435 27489 8447 27523
rect 8389 27483 8447 27489
rect 9306 27480 9312 27532
rect 9364 27520 9370 27532
rect 10229 27523 10287 27529
rect 10229 27520 10241 27523
rect 9364 27492 10241 27520
rect 9364 27480 9370 27492
rect 10229 27489 10241 27492
rect 10275 27489 10287 27523
rect 10229 27483 10287 27489
rect 11054 27480 11060 27532
rect 11112 27520 11118 27532
rect 12158 27520 12164 27532
rect 11112 27492 12164 27520
rect 11112 27480 11118 27492
rect 12158 27480 12164 27492
rect 12216 27520 12222 27532
rect 12253 27523 12311 27529
rect 12253 27520 12265 27523
rect 12216 27492 12265 27520
rect 12216 27480 12222 27492
rect 12253 27489 12265 27492
rect 12299 27520 12311 27523
rect 12342 27520 12348 27532
rect 12299 27492 12348 27520
rect 12299 27489 12311 27492
rect 12253 27483 12311 27489
rect 12342 27480 12348 27492
rect 12400 27480 12406 27532
rect 12526 27480 12532 27532
rect 12584 27520 12590 27532
rect 15856 27529 15884 27560
rect 18506 27548 18512 27600
rect 18564 27588 18570 27600
rect 18877 27591 18935 27597
rect 18877 27588 18889 27591
rect 18564 27560 18889 27588
rect 18564 27548 18570 27560
rect 18877 27557 18889 27560
rect 18923 27557 18935 27591
rect 20438 27588 20444 27600
rect 18877 27551 18935 27557
rect 19904 27560 20444 27588
rect 13265 27523 13323 27529
rect 13265 27520 13277 27523
rect 12584 27492 13277 27520
rect 12584 27480 12590 27492
rect 13265 27489 13277 27492
rect 13311 27489 13323 27523
rect 13265 27483 13323 27489
rect 15841 27523 15899 27529
rect 15841 27489 15853 27523
rect 15887 27489 15899 27523
rect 18230 27520 18236 27532
rect 18143 27492 18236 27520
rect 15841 27483 15899 27489
rect 18230 27480 18236 27492
rect 18288 27480 18294 27532
rect 18414 27520 18420 27532
rect 18375 27492 18420 27520
rect 18414 27480 18420 27492
rect 18472 27520 18478 27532
rect 19904 27529 19932 27560
rect 20438 27548 20444 27560
rect 20496 27548 20502 27600
rect 20806 27588 20812 27600
rect 20548 27560 20812 27588
rect 19889 27523 19947 27529
rect 19889 27520 19901 27523
rect 18472 27492 19901 27520
rect 18472 27480 18478 27492
rect 19889 27489 19901 27492
rect 19935 27489 19947 27523
rect 19889 27483 19947 27489
rect 20073 27523 20131 27529
rect 20073 27489 20085 27523
rect 20119 27520 20131 27523
rect 20548 27520 20576 27560
rect 20806 27548 20812 27560
rect 20864 27548 20870 27600
rect 23474 27588 23480 27600
rect 23435 27560 23480 27588
rect 23474 27548 23480 27560
rect 23532 27548 23538 27600
rect 22833 27523 22891 27529
rect 20119 27492 20576 27520
rect 20732 27492 22094 27520
rect 20119 27489 20131 27492
rect 20073 27483 20131 27489
rect 7377 27455 7435 27461
rect 7377 27421 7389 27455
rect 7423 27452 7435 27455
rect 8754 27452 8760 27464
rect 7423 27424 8760 27452
rect 7423 27421 7435 27424
rect 7377 27415 7435 27421
rect 8754 27412 8760 27424
rect 8812 27412 8818 27464
rect 9582 27452 9588 27464
rect 9543 27424 9588 27452
rect 9582 27412 9588 27424
rect 9640 27412 9646 27464
rect 14550 27452 14556 27464
rect 14511 27424 14556 27452
rect 14550 27412 14556 27424
rect 14608 27412 14614 27464
rect 15197 27455 15255 27461
rect 15197 27421 15209 27455
rect 15243 27421 15255 27455
rect 18248 27452 18276 27480
rect 19334 27452 19340 27464
rect 18248 27424 19340 27452
rect 15197 27415 15255 27421
rect 8205 27387 8263 27393
rect 8205 27353 8217 27387
rect 8251 27384 8263 27387
rect 9674 27384 9680 27396
rect 8251 27356 9680 27384
rect 8251 27353 8263 27356
rect 8205 27347 8263 27353
rect 9674 27344 9680 27356
rect 9732 27344 9738 27396
rect 10505 27387 10563 27393
rect 10505 27384 10517 27387
rect 9784 27356 10517 27384
rect 7837 27319 7895 27325
rect 7837 27285 7849 27319
rect 7883 27316 7895 27319
rect 7926 27316 7932 27328
rect 7883 27288 7932 27316
rect 7883 27285 7895 27288
rect 7837 27279 7895 27285
rect 7926 27276 7932 27288
rect 7984 27276 7990 27328
rect 8297 27319 8355 27325
rect 8297 27285 8309 27319
rect 8343 27316 8355 27319
rect 9214 27316 9220 27328
rect 8343 27288 9220 27316
rect 8343 27285 8355 27288
rect 8297 27279 8355 27285
rect 9214 27276 9220 27288
rect 9272 27276 9278 27328
rect 9784 27325 9812 27356
rect 10505 27353 10517 27356
rect 10551 27353 10563 27387
rect 11790 27384 11796 27396
rect 11730 27356 11796 27384
rect 10505 27347 10563 27353
rect 11790 27344 11796 27356
rect 11848 27344 11854 27396
rect 12342 27344 12348 27396
rect 12400 27384 12406 27396
rect 13173 27387 13231 27393
rect 13173 27384 13185 27387
rect 12400 27356 13185 27384
rect 12400 27344 12406 27356
rect 13173 27353 13185 27356
rect 13219 27353 13231 27387
rect 13173 27347 13231 27353
rect 13722 27344 13728 27396
rect 13780 27384 13786 27396
rect 15212 27384 15240 27415
rect 19334 27412 19340 27424
rect 19392 27412 19398 27464
rect 19797 27455 19855 27461
rect 19797 27421 19809 27455
rect 19843 27452 19855 27455
rect 20732 27452 20760 27492
rect 19843 27424 20760 27452
rect 20809 27455 20867 27461
rect 19843 27421 19855 27424
rect 19797 27415 19855 27421
rect 20809 27421 20821 27455
rect 20855 27421 20867 27455
rect 21266 27452 21272 27464
rect 21227 27424 21272 27452
rect 20809 27415 20867 27421
rect 13780 27356 15240 27384
rect 13780 27344 13786 27356
rect 9769 27319 9827 27325
rect 9769 27285 9781 27319
rect 9815 27285 9827 27319
rect 9769 27279 9827 27285
rect 11146 27276 11152 27328
rect 11204 27316 11210 27328
rect 12713 27319 12771 27325
rect 12713 27316 12725 27319
rect 11204 27288 12725 27316
rect 11204 27276 11210 27288
rect 12713 27285 12725 27288
rect 12759 27285 12771 27319
rect 13078 27316 13084 27328
rect 13039 27288 13084 27316
rect 12713 27279 12771 27285
rect 13078 27276 13084 27288
rect 13136 27276 13142 27328
rect 14182 27276 14188 27328
rect 14240 27316 14246 27328
rect 14369 27319 14427 27325
rect 14369 27316 14381 27319
rect 14240 27288 14381 27316
rect 14240 27276 14246 27288
rect 14369 27285 14381 27288
rect 14415 27285 14427 27319
rect 15212 27316 15240 27356
rect 15289 27387 15347 27393
rect 15289 27353 15301 27387
rect 15335 27384 15347 27387
rect 15335 27356 16606 27384
rect 15335 27353 15347 27356
rect 15289 27347 15347 27353
rect 18874 27344 18880 27396
rect 18932 27384 18938 27396
rect 20824 27384 20852 27415
rect 21266 27412 21272 27424
rect 21324 27412 21330 27464
rect 18932 27356 20852 27384
rect 22066 27384 22094 27492
rect 22833 27489 22845 27523
rect 22879 27520 22891 27523
rect 22879 27492 23520 27520
rect 22879 27489 22891 27492
rect 22833 27483 22891 27489
rect 23492 27464 23520 27492
rect 22557 27455 22615 27461
rect 22557 27421 22569 27455
rect 22603 27452 22615 27455
rect 23198 27452 23204 27464
rect 22603 27424 23204 27452
rect 22603 27421 22615 27424
rect 22557 27415 22615 27421
rect 23198 27412 23204 27424
rect 23256 27412 23262 27464
rect 23474 27412 23480 27464
rect 23532 27412 23538 27464
rect 23584 27461 23612 27628
rect 28810 27616 28816 27668
rect 28868 27656 28874 27668
rect 28905 27659 28963 27665
rect 28905 27656 28917 27659
rect 28868 27628 28917 27656
rect 28868 27616 28874 27628
rect 28905 27625 28917 27628
rect 28951 27625 28963 27659
rect 28905 27619 28963 27625
rect 35434 27616 35440 27668
rect 35492 27656 35498 27668
rect 35621 27659 35679 27665
rect 35621 27656 35633 27659
rect 35492 27628 35633 27656
rect 35492 27616 35498 27628
rect 35621 27625 35633 27628
rect 35667 27625 35679 27659
rect 35621 27619 35679 27625
rect 31573 27591 31631 27597
rect 31573 27557 31585 27591
rect 31619 27588 31631 27591
rect 31754 27588 31760 27600
rect 31619 27560 31760 27588
rect 31619 27557 31631 27560
rect 31573 27551 31631 27557
rect 31754 27548 31760 27560
rect 31812 27548 31818 27600
rect 34606 27588 34612 27600
rect 32324 27560 34612 27588
rect 23658 27480 23664 27532
rect 23716 27520 23722 27532
rect 24854 27520 24860 27532
rect 23716 27492 24860 27520
rect 23716 27480 23722 27492
rect 24854 27480 24860 27492
rect 24912 27520 24918 27532
rect 24949 27523 25007 27529
rect 24949 27520 24961 27523
rect 24912 27492 24961 27520
rect 24912 27480 24918 27492
rect 24949 27489 24961 27492
rect 24995 27520 25007 27523
rect 30469 27523 30527 27529
rect 24995 27492 27200 27520
rect 24995 27489 25007 27492
rect 24949 27483 25007 27489
rect 27172 27464 27200 27492
rect 30469 27489 30481 27523
rect 30515 27520 30527 27523
rect 32324 27520 32352 27560
rect 34606 27548 34612 27560
rect 34664 27548 34670 27600
rect 36170 27588 36176 27600
rect 36131 27560 36176 27588
rect 36170 27548 36176 27560
rect 36228 27548 36234 27600
rect 37090 27588 37096 27600
rect 37051 27560 37096 27588
rect 37090 27548 37096 27560
rect 37148 27548 37154 27600
rect 32490 27520 32496 27532
rect 30515 27492 32352 27520
rect 32451 27492 32496 27520
rect 30515 27489 30527 27492
rect 30469 27483 30527 27489
rect 32490 27480 32496 27492
rect 32548 27480 32554 27532
rect 33318 27480 33324 27532
rect 33376 27520 33382 27532
rect 33413 27523 33471 27529
rect 33413 27520 33425 27523
rect 33376 27492 33425 27520
rect 33376 27480 33382 27492
rect 33413 27489 33425 27492
rect 33459 27489 33471 27523
rect 33413 27483 33471 27489
rect 33873 27523 33931 27529
rect 33873 27489 33885 27523
rect 33919 27489 33931 27523
rect 33873 27483 33931 27489
rect 23569 27455 23627 27461
rect 23569 27421 23581 27455
rect 23615 27452 23627 27455
rect 24670 27452 24676 27464
rect 23615 27424 24676 27452
rect 23615 27421 23627 27424
rect 23569 27415 23627 27421
rect 24670 27412 24676 27424
rect 24728 27412 24734 27464
rect 27154 27452 27160 27464
rect 27115 27424 27160 27452
rect 27154 27412 27160 27424
rect 27212 27412 27218 27464
rect 30377 27455 30435 27461
rect 30377 27421 30389 27455
rect 30423 27421 30435 27455
rect 30377 27415 30435 27421
rect 24946 27384 24952 27396
rect 22066 27356 24952 27384
rect 18932 27344 18938 27356
rect 24946 27344 24952 27356
rect 25004 27344 25010 27396
rect 25222 27384 25228 27396
rect 25183 27356 25228 27384
rect 25222 27344 25228 27356
rect 25280 27344 25286 27396
rect 26878 27384 26884 27396
rect 26450 27356 26884 27384
rect 26878 27344 26884 27356
rect 26936 27344 26942 27396
rect 27430 27384 27436 27396
rect 27391 27356 27436 27384
rect 27430 27344 27436 27356
rect 27488 27344 27494 27396
rect 27522 27344 27528 27396
rect 27580 27384 27586 27396
rect 30392 27384 30420 27415
rect 31018 27412 31024 27464
rect 31076 27452 31082 27464
rect 31205 27455 31263 27461
rect 31205 27452 31217 27455
rect 31076 27424 31217 27452
rect 31076 27412 31082 27424
rect 31205 27421 31217 27424
rect 31251 27421 31263 27455
rect 31386 27452 31392 27464
rect 31347 27424 31392 27452
rect 31205 27415 31263 27421
rect 31386 27412 31392 27424
rect 31444 27412 31450 27464
rect 32401 27455 32459 27461
rect 32401 27421 32413 27455
rect 32447 27452 32459 27455
rect 32858 27452 32864 27464
rect 32447 27424 32864 27452
rect 32447 27421 32459 27424
rect 32401 27415 32459 27421
rect 31570 27384 31576 27396
rect 27580 27356 27922 27384
rect 30392 27356 31576 27384
rect 27580 27344 27586 27356
rect 31570 27344 31576 27356
rect 31628 27344 31634 27396
rect 16482 27316 16488 27328
rect 15212 27288 16488 27316
rect 14369 27279 14427 27285
rect 16482 27276 16488 27288
rect 16540 27276 16546 27328
rect 17586 27316 17592 27328
rect 17547 27288 17592 27316
rect 17586 27276 17592 27288
rect 17644 27276 17650 27328
rect 18414 27276 18420 27328
rect 18472 27316 18478 27328
rect 18509 27319 18567 27325
rect 18509 27316 18521 27319
rect 18472 27288 18521 27316
rect 18472 27276 18478 27288
rect 18509 27285 18521 27288
rect 18555 27285 18567 27319
rect 19426 27316 19432 27328
rect 19387 27288 19432 27316
rect 18509 27279 18567 27285
rect 19426 27276 19432 27288
rect 19484 27276 19490 27328
rect 20622 27316 20628 27328
rect 20583 27288 20628 27316
rect 20622 27276 20628 27288
rect 20680 27276 20686 27328
rect 21358 27316 21364 27328
rect 21319 27288 21364 27316
rect 21358 27276 21364 27288
rect 21416 27276 21422 27328
rect 22186 27316 22192 27328
rect 22147 27288 22192 27316
rect 22186 27276 22192 27288
rect 22244 27276 22250 27328
rect 22646 27316 22652 27328
rect 22607 27288 22652 27316
rect 22646 27276 22652 27288
rect 22704 27276 22710 27328
rect 24578 27276 24584 27328
rect 24636 27316 24642 27328
rect 26697 27319 26755 27325
rect 26697 27316 26709 27319
rect 24636 27288 26709 27316
rect 24636 27276 24642 27288
rect 26697 27285 26709 27288
rect 26743 27316 26755 27319
rect 28350 27316 28356 27328
rect 26743 27288 28356 27316
rect 26743 27285 26755 27288
rect 26697 27279 26755 27285
rect 28350 27276 28356 27288
rect 28408 27276 28414 27328
rect 30742 27316 30748 27328
rect 30703 27288 30748 27316
rect 30742 27276 30748 27288
rect 30800 27276 30806 27328
rect 30834 27276 30840 27328
rect 30892 27316 30898 27328
rect 32416 27316 32444 27415
rect 32858 27412 32864 27424
rect 32916 27412 32922 27464
rect 33505 27455 33563 27461
rect 33505 27421 33517 27455
rect 33551 27421 33563 27455
rect 33888 27452 33916 27483
rect 34790 27480 34796 27532
rect 34848 27520 34854 27532
rect 34977 27523 35035 27529
rect 34977 27520 34989 27523
rect 34848 27492 34989 27520
rect 34848 27480 34854 27492
rect 34977 27489 34989 27492
rect 35023 27489 35035 27523
rect 34977 27483 35035 27489
rect 35158 27480 35164 27532
rect 35216 27520 35222 27532
rect 36630 27520 36636 27532
rect 35216 27492 36636 27520
rect 35216 27480 35222 27492
rect 36630 27480 36636 27492
rect 36688 27480 36694 27532
rect 35253 27455 35311 27461
rect 35253 27452 35265 27455
rect 33888 27424 35265 27452
rect 33505 27415 33563 27421
rect 35253 27421 35265 27424
rect 35299 27421 35311 27455
rect 35253 27415 35311 27421
rect 36265 27455 36323 27461
rect 36265 27421 36277 27455
rect 36311 27452 36323 27455
rect 36354 27452 36360 27464
rect 36311 27424 36360 27452
rect 36311 27421 36323 27424
rect 36265 27415 36323 27421
rect 33042 27384 33048 27396
rect 32784 27356 33048 27384
rect 32784 27325 32812 27356
rect 33042 27344 33048 27356
rect 33100 27384 33106 27396
rect 33520 27384 33548 27415
rect 36354 27412 36360 27424
rect 36412 27412 36418 27464
rect 36909 27455 36967 27461
rect 36909 27421 36921 27455
rect 36955 27452 36967 27455
rect 36998 27452 37004 27464
rect 36955 27424 37004 27452
rect 36955 27421 36967 27424
rect 36909 27415 36967 27421
rect 36998 27412 37004 27424
rect 37056 27412 37062 27464
rect 33100 27356 35296 27384
rect 33100 27344 33106 27356
rect 30892 27288 32444 27316
rect 32769 27319 32827 27325
rect 30892 27276 30898 27288
rect 32769 27285 32781 27319
rect 32815 27285 32827 27319
rect 32769 27279 32827 27285
rect 32858 27276 32864 27328
rect 32916 27316 32922 27328
rect 35158 27316 35164 27328
rect 32916 27288 35164 27316
rect 32916 27276 32922 27288
rect 35158 27276 35164 27288
rect 35216 27276 35222 27328
rect 35268 27316 35296 27356
rect 36446 27316 36452 27328
rect 35268 27288 36452 27316
rect 36446 27276 36452 27288
rect 36504 27276 36510 27328
rect 1104 27226 37628 27248
rect 1104 27174 4874 27226
rect 4926 27174 4938 27226
rect 4990 27174 5002 27226
rect 5054 27174 5066 27226
rect 5118 27174 5130 27226
rect 5182 27174 35594 27226
rect 35646 27174 35658 27226
rect 35710 27174 35722 27226
rect 35774 27174 35786 27226
rect 35838 27174 35850 27226
rect 35902 27174 37628 27226
rect 1104 27152 37628 27174
rect 9125 27115 9183 27121
rect 9125 27081 9137 27115
rect 9171 27112 9183 27115
rect 9214 27112 9220 27124
rect 9171 27084 9220 27112
rect 9171 27081 9183 27084
rect 9125 27075 9183 27081
rect 9214 27072 9220 27084
rect 9272 27072 9278 27124
rect 9582 27112 9588 27124
rect 9543 27084 9588 27112
rect 9582 27072 9588 27084
rect 9640 27072 9646 27124
rect 9674 27072 9680 27124
rect 9732 27112 9738 27124
rect 11701 27115 11759 27121
rect 11701 27112 11713 27115
rect 9732 27084 11713 27112
rect 9732 27072 9738 27084
rect 11701 27081 11713 27084
rect 11747 27081 11759 27115
rect 12158 27112 12164 27124
rect 12119 27084 12164 27112
rect 11701 27075 11759 27081
rect 12158 27072 12164 27084
rect 12216 27072 12222 27124
rect 13722 27112 13728 27124
rect 13280 27084 13728 27112
rect 8386 27004 8392 27056
rect 8444 27004 8450 27056
rect 9232 27044 9260 27072
rect 10045 27047 10103 27053
rect 10045 27044 10057 27047
rect 9232 27016 10057 27044
rect 10045 27013 10057 27016
rect 10091 27013 10103 27047
rect 10045 27007 10103 27013
rect 11238 27004 11244 27056
rect 11296 27044 11302 27056
rect 12069 27047 12127 27053
rect 12069 27044 12081 27047
rect 11296 27016 12081 27044
rect 11296 27004 11302 27016
rect 12069 27013 12081 27016
rect 12115 27044 12127 27047
rect 12342 27044 12348 27056
rect 12115 27016 12348 27044
rect 12115 27013 12127 27016
rect 12069 27007 12127 27013
rect 12342 27004 12348 27016
rect 12400 27004 12406 27056
rect 9953 26979 10011 26985
rect 9953 26945 9965 26979
rect 9999 26976 10011 26979
rect 11054 26976 11060 26988
rect 9999 26948 11060 26976
rect 9999 26945 10011 26948
rect 9953 26939 10011 26945
rect 11054 26936 11060 26948
rect 11112 26936 11118 26988
rect 11149 26979 11207 26985
rect 11149 26945 11161 26979
rect 11195 26976 11207 26979
rect 11698 26976 11704 26988
rect 11195 26948 11704 26976
rect 11195 26945 11207 26948
rect 11149 26939 11207 26945
rect 11698 26936 11704 26948
rect 11756 26976 11762 26988
rect 13280 26976 13308 27084
rect 13722 27072 13728 27084
rect 13780 27072 13786 27124
rect 14550 27072 14556 27124
rect 14608 27112 14614 27124
rect 15473 27115 15531 27121
rect 15473 27112 15485 27115
rect 14608 27084 15485 27112
rect 14608 27072 14614 27084
rect 15473 27081 15485 27084
rect 15519 27081 15531 27115
rect 21358 27112 21364 27124
rect 15473 27075 15531 27081
rect 19352 27084 21364 27112
rect 13538 27044 13544 27056
rect 13499 27016 13544 27044
rect 13538 27004 13544 27016
rect 13596 27004 13602 27056
rect 13630 27004 13636 27056
rect 13688 27044 13694 27056
rect 13688 27016 14030 27044
rect 13688 27004 13694 27016
rect 16758 27004 16764 27056
rect 16816 27044 16822 27056
rect 19352 27044 19380 27084
rect 21358 27072 21364 27084
rect 21416 27072 21422 27124
rect 22646 27072 22652 27124
rect 22704 27112 22710 27124
rect 24210 27112 24216 27124
rect 22704 27084 24216 27112
rect 22704 27072 22710 27084
rect 24210 27072 24216 27084
rect 24268 27112 24274 27124
rect 24673 27115 24731 27121
rect 24673 27112 24685 27115
rect 24268 27084 24685 27112
rect 24268 27072 24274 27084
rect 24673 27081 24685 27084
rect 24719 27081 24731 27115
rect 24673 27075 24731 27081
rect 25133 27115 25191 27121
rect 25133 27081 25145 27115
rect 25179 27081 25191 27115
rect 25133 27075 25191 27081
rect 16816 27016 17080 27044
rect 18998 27016 19380 27044
rect 19429 27047 19487 27053
rect 16816 27004 16822 27016
rect 17052 26985 17080 27016
rect 19429 27013 19441 27047
rect 19475 27044 19487 27047
rect 20622 27044 20628 27056
rect 19475 27016 20628 27044
rect 19475 27013 19487 27016
rect 19429 27007 19487 27013
rect 20622 27004 20628 27016
rect 20680 27004 20686 27056
rect 22833 27047 22891 27053
rect 22833 27044 22845 27047
rect 22066 27016 22845 27044
rect 11756 26948 13308 26976
rect 15841 26979 15899 26985
rect 11756 26936 11762 26948
rect 15841 26945 15853 26979
rect 15887 26976 15899 26979
rect 17037 26979 17095 26985
rect 15887 26948 16988 26976
rect 15887 26945 15899 26948
rect 15841 26939 15899 26945
rect 7377 26911 7435 26917
rect 7377 26877 7389 26911
rect 7423 26877 7435 26911
rect 7377 26871 7435 26877
rect 7653 26911 7711 26917
rect 7653 26877 7665 26911
rect 7699 26908 7711 26911
rect 7742 26908 7748 26920
rect 7699 26880 7748 26908
rect 7699 26877 7711 26880
rect 7653 26871 7711 26877
rect 7392 26772 7420 26871
rect 7742 26868 7748 26880
rect 7800 26868 7806 26920
rect 10229 26911 10287 26917
rect 10229 26877 10241 26911
rect 10275 26908 10287 26911
rect 12345 26911 12403 26917
rect 10275 26880 11744 26908
rect 10275 26877 10287 26880
rect 10229 26871 10287 26877
rect 9030 26772 9036 26784
rect 7392 26744 9036 26772
rect 9030 26732 9036 26744
rect 9088 26732 9094 26784
rect 11057 26775 11115 26781
rect 11057 26741 11069 26775
rect 11103 26772 11115 26775
rect 11422 26772 11428 26784
rect 11103 26744 11428 26772
rect 11103 26741 11115 26744
rect 11057 26735 11115 26741
rect 11422 26732 11428 26744
rect 11480 26732 11486 26784
rect 11716 26772 11744 26880
rect 12345 26877 12357 26911
rect 12391 26908 12403 26911
rect 12710 26908 12716 26920
rect 12391 26880 12716 26908
rect 12391 26877 12403 26880
rect 12345 26871 12403 26877
rect 12710 26868 12716 26880
rect 12768 26868 12774 26920
rect 13265 26911 13323 26917
rect 13265 26877 13277 26911
rect 13311 26877 13323 26911
rect 15010 26908 15016 26920
rect 14971 26880 15016 26908
rect 13265 26871 13323 26877
rect 11790 26800 11796 26852
rect 11848 26840 11854 26852
rect 13280 26840 13308 26871
rect 15010 26868 15016 26880
rect 15068 26908 15074 26920
rect 15933 26911 15991 26917
rect 15933 26908 15945 26911
rect 15068 26880 15945 26908
rect 15068 26868 15074 26880
rect 15933 26877 15945 26880
rect 15979 26877 15991 26911
rect 15933 26871 15991 26877
rect 16117 26911 16175 26917
rect 16117 26877 16129 26911
rect 16163 26877 16175 26911
rect 16960 26908 16988 26948
rect 17037 26945 17049 26979
rect 17083 26945 17095 26979
rect 17037 26939 17095 26945
rect 20070 26936 20076 26988
rect 20128 26976 20134 26988
rect 20257 26979 20315 26985
rect 20257 26976 20269 26979
rect 20128 26948 20269 26976
rect 20128 26936 20134 26948
rect 20257 26945 20269 26948
rect 20303 26976 20315 26979
rect 20714 26976 20720 26988
rect 20303 26948 20720 26976
rect 20303 26945 20315 26948
rect 20257 26939 20315 26945
rect 20714 26936 20720 26948
rect 20772 26976 20778 26988
rect 22066 26976 22094 27016
rect 22833 27013 22845 27016
rect 22879 27013 22891 27047
rect 23658 27044 23664 27056
rect 23619 27016 23664 27044
rect 22833 27007 22891 27013
rect 23658 27004 23664 27016
rect 23716 27004 23722 27056
rect 24578 27004 24584 27056
rect 24636 27044 24642 27056
rect 24765 27047 24823 27053
rect 24765 27044 24777 27047
rect 24636 27016 24777 27044
rect 24636 27004 24642 27016
rect 24765 27013 24777 27016
rect 24811 27013 24823 27047
rect 24765 27007 24823 27013
rect 20772 26948 22094 26976
rect 20772 26936 20778 26948
rect 22186 26936 22192 26988
rect 22244 26976 22250 26988
rect 25148 26976 25176 27075
rect 25222 27072 25228 27124
rect 25280 27112 25286 27124
rect 25593 27115 25651 27121
rect 25593 27112 25605 27115
rect 25280 27084 25605 27112
rect 25280 27072 25286 27084
rect 25593 27081 25605 27084
rect 25639 27081 25651 27115
rect 25593 27075 25651 27081
rect 26421 27115 26479 27121
rect 26421 27081 26433 27115
rect 26467 27112 26479 27115
rect 27430 27112 27436 27124
rect 26467 27084 27436 27112
rect 26467 27081 26479 27084
rect 26421 27075 26479 27081
rect 27430 27072 27436 27084
rect 27488 27072 27494 27124
rect 28721 27115 28779 27121
rect 28721 27081 28733 27115
rect 28767 27112 28779 27115
rect 29178 27112 29184 27124
rect 28767 27084 29184 27112
rect 28767 27081 28779 27084
rect 28721 27075 28779 27081
rect 29178 27072 29184 27084
rect 29236 27072 29242 27124
rect 30742 27112 30748 27124
rect 30703 27084 30748 27112
rect 30742 27072 30748 27084
rect 30800 27072 30806 27124
rect 32950 27112 32956 27124
rect 30852 27084 32956 27112
rect 28626 27004 28632 27056
rect 28684 27044 28690 27056
rect 30852 27044 30880 27084
rect 32950 27072 32956 27084
rect 33008 27072 33014 27124
rect 33318 27072 33324 27124
rect 33376 27112 33382 27124
rect 33376 27084 36676 27112
rect 33376 27072 33382 27084
rect 31386 27044 31392 27056
rect 28684 27016 30880 27044
rect 30944 27016 31392 27044
rect 28684 27004 28690 27016
rect 25777 26979 25835 26985
rect 25777 26976 25789 26979
rect 22244 26948 22289 26976
rect 25148 26948 25789 26976
rect 22244 26936 22250 26948
rect 25777 26945 25789 26948
rect 25823 26945 25835 26979
rect 25777 26939 25835 26945
rect 26142 26936 26148 26988
rect 26200 26976 26206 26988
rect 26237 26979 26295 26985
rect 26237 26976 26249 26979
rect 26200 26948 26249 26976
rect 26200 26936 26206 26948
rect 26237 26945 26249 26948
rect 26283 26945 26295 26979
rect 26237 26939 26295 26945
rect 26694 26936 26700 26988
rect 26752 26976 26758 26988
rect 27157 26979 27215 26985
rect 27157 26976 27169 26979
rect 26752 26948 27169 26976
rect 26752 26936 26758 26948
rect 27157 26945 27169 26948
rect 27203 26945 27215 26979
rect 28350 26976 28356 26988
rect 28311 26948 28356 26976
rect 27157 26939 27215 26945
rect 28350 26936 28356 26948
rect 28408 26936 28414 26988
rect 28534 26976 28540 26988
rect 28495 26948 28540 26976
rect 28534 26936 28540 26948
rect 28592 26936 28598 26988
rect 29181 26979 29239 26985
rect 29181 26945 29193 26979
rect 29227 26945 29239 26979
rect 29181 26939 29239 26945
rect 18966 26908 18972 26920
rect 16960 26880 18972 26908
rect 16117 26871 16175 26877
rect 11848 26812 13308 26840
rect 11848 26800 11854 26812
rect 15102 26800 15108 26852
rect 15160 26840 15166 26852
rect 16132 26840 16160 26871
rect 18966 26868 18972 26880
rect 19024 26868 19030 26920
rect 19702 26908 19708 26920
rect 19663 26880 19708 26908
rect 19702 26868 19708 26880
rect 19760 26908 19766 26920
rect 20993 26911 21051 26917
rect 20993 26908 21005 26911
rect 19760 26880 21005 26908
rect 19760 26868 19766 26880
rect 20993 26877 21005 26880
rect 21039 26877 21051 26911
rect 24581 26911 24639 26917
rect 20993 26871 21051 26877
rect 21100 26880 22094 26908
rect 17402 26840 17408 26852
rect 15160 26812 17408 26840
rect 15160 26800 15166 26812
rect 17402 26800 17408 26812
rect 17460 26800 17466 26852
rect 19794 26800 19800 26852
rect 19852 26840 19858 26852
rect 21100 26840 21128 26880
rect 19852 26812 21128 26840
rect 22066 26840 22094 26880
rect 24581 26877 24593 26911
rect 24627 26908 24639 26911
rect 25130 26908 25136 26920
rect 24627 26880 25136 26908
rect 24627 26877 24639 26880
rect 24581 26871 24639 26877
rect 25130 26868 25136 26880
rect 25188 26868 25194 26920
rect 26602 26868 26608 26920
rect 26660 26908 26666 26920
rect 27338 26908 27344 26920
rect 26660 26880 27344 26908
rect 26660 26868 26666 26880
rect 27338 26868 27344 26880
rect 27396 26908 27402 26920
rect 29196 26908 29224 26939
rect 30466 26936 30472 26988
rect 30524 26976 30530 26988
rect 30653 26979 30711 26985
rect 30653 26976 30665 26979
rect 30524 26948 30665 26976
rect 30524 26936 30530 26948
rect 30653 26945 30665 26948
rect 30699 26976 30711 26979
rect 30944 26976 30972 27016
rect 31386 27004 31392 27016
rect 31444 27044 31450 27056
rect 33413 27047 33471 27053
rect 31444 27016 33364 27044
rect 31444 27004 31450 27016
rect 31573 26979 31631 26985
rect 31573 26976 31585 26979
rect 30699 26948 30972 26976
rect 31128 26948 31585 26976
rect 30699 26945 30711 26948
rect 30653 26939 30711 26945
rect 30558 26908 30564 26920
rect 27396 26880 29224 26908
rect 30519 26880 30564 26908
rect 27396 26868 27402 26880
rect 30558 26868 30564 26880
rect 30616 26868 30622 26920
rect 28534 26840 28540 26852
rect 22066 26812 28540 26840
rect 19852 26800 19858 26812
rect 28534 26800 28540 26812
rect 28592 26840 28598 26852
rect 30834 26840 30840 26852
rect 28592 26812 30840 26840
rect 28592 26800 28598 26812
rect 30834 26800 30840 26812
rect 30892 26800 30898 26852
rect 31128 26849 31156 26948
rect 31573 26945 31585 26948
rect 31619 26945 31631 26979
rect 31573 26939 31631 26945
rect 32306 26936 32312 26988
rect 32364 26976 32370 26988
rect 33336 26985 33364 27016
rect 33413 27013 33425 27047
rect 33459 27044 33471 27047
rect 33502 27044 33508 27056
rect 33459 27016 33508 27044
rect 33459 27013 33471 27016
rect 33413 27007 33471 27013
rect 33502 27004 33508 27016
rect 33560 27004 33566 27056
rect 34164 27016 35848 27044
rect 32493 26979 32551 26985
rect 32493 26976 32505 26979
rect 32364 26948 32505 26976
rect 32364 26936 32370 26948
rect 32493 26945 32505 26948
rect 32539 26945 32551 26979
rect 32493 26939 32551 26945
rect 33321 26979 33379 26985
rect 33321 26945 33333 26979
rect 33367 26945 33379 26979
rect 34164 26976 34192 27016
rect 35820 26988 35848 27016
rect 33321 26939 33379 26945
rect 33428 26948 34192 26976
rect 32401 26911 32459 26917
rect 32401 26877 32413 26911
rect 32447 26908 32459 26911
rect 32447 26880 32536 26908
rect 32447 26877 32459 26880
rect 32401 26871 32459 26877
rect 32508 26852 32536 26880
rect 32950 26868 32956 26920
rect 33008 26908 33014 26920
rect 33428 26908 33456 26948
rect 34238 26936 34244 26988
rect 34296 26976 34302 26988
rect 34609 26979 34667 26985
rect 34609 26976 34621 26979
rect 34296 26948 34621 26976
rect 34296 26936 34302 26948
rect 34609 26945 34621 26948
rect 34655 26945 34667 26979
rect 35802 26976 35808 26988
rect 35715 26948 35808 26976
rect 34609 26939 34667 26945
rect 35802 26936 35808 26948
rect 35860 26936 35866 26988
rect 36446 26976 36452 26988
rect 36407 26948 36452 26976
rect 36446 26936 36452 26948
rect 36504 26936 36510 26988
rect 36648 26985 36676 27084
rect 36633 26979 36691 26985
rect 36633 26945 36645 26979
rect 36679 26945 36691 26979
rect 36633 26939 36691 26945
rect 33008 26880 33456 26908
rect 34425 26911 34483 26917
rect 33008 26868 33014 26880
rect 34425 26877 34437 26911
rect 34471 26877 34483 26911
rect 34425 26871 34483 26877
rect 34517 26911 34575 26917
rect 34517 26877 34529 26911
rect 34563 26877 34575 26911
rect 34517 26871 34575 26877
rect 31113 26843 31171 26849
rect 31113 26809 31125 26843
rect 31159 26809 31171 26843
rect 31113 26803 31171 26809
rect 32490 26800 32496 26852
rect 32548 26800 32554 26852
rect 12526 26772 12532 26784
rect 11716 26744 12532 26772
rect 12526 26732 12532 26744
rect 12584 26732 12590 26784
rect 17129 26775 17187 26781
rect 17129 26741 17141 26775
rect 17175 26772 17187 26775
rect 17218 26772 17224 26784
rect 17175 26744 17224 26772
rect 17175 26741 17187 26744
rect 17129 26735 17187 26741
rect 17218 26732 17224 26744
rect 17276 26732 17282 26784
rect 17957 26775 18015 26781
rect 17957 26741 17969 26775
rect 18003 26772 18015 26775
rect 18414 26772 18420 26784
rect 18003 26744 18420 26772
rect 18003 26741 18015 26744
rect 17957 26735 18015 26741
rect 18414 26732 18420 26744
rect 18472 26732 18478 26784
rect 19610 26732 19616 26784
rect 19668 26772 19674 26784
rect 19886 26772 19892 26784
rect 19668 26744 19892 26772
rect 19668 26732 19674 26744
rect 19886 26732 19892 26744
rect 19944 26732 19950 26784
rect 20990 26732 20996 26784
rect 21048 26772 21054 26784
rect 22005 26775 22063 26781
rect 22005 26772 22017 26775
rect 21048 26744 22017 26772
rect 21048 26732 21054 26744
rect 22005 26741 22017 26744
rect 22051 26741 22063 26775
rect 22005 26735 22063 26741
rect 22370 26732 22376 26784
rect 22428 26772 22434 26784
rect 28442 26772 28448 26784
rect 22428 26744 28448 26772
rect 22428 26732 22434 26744
rect 28442 26732 28448 26744
rect 28500 26732 28506 26784
rect 29270 26772 29276 26784
rect 29231 26744 29276 26772
rect 29270 26732 29276 26744
rect 29328 26732 29334 26784
rect 31662 26732 31668 26784
rect 31720 26772 31726 26784
rect 31757 26775 31815 26781
rect 31757 26772 31769 26775
rect 31720 26744 31769 26772
rect 31720 26732 31726 26744
rect 31757 26741 31769 26744
rect 31803 26741 31815 26775
rect 31757 26735 31815 26741
rect 32769 26775 32827 26781
rect 32769 26741 32781 26775
rect 32815 26772 32827 26775
rect 32950 26772 32956 26784
rect 32815 26744 32956 26772
rect 32815 26741 32827 26744
rect 32769 26735 32827 26741
rect 32950 26732 32956 26744
rect 33008 26772 33014 26784
rect 33962 26772 33968 26784
rect 33008 26744 33968 26772
rect 33008 26732 33014 26744
rect 33962 26732 33968 26744
rect 34020 26732 34026 26784
rect 34440 26772 34468 26871
rect 34532 26840 34560 26871
rect 34790 26868 34796 26920
rect 34848 26908 34854 26920
rect 35713 26911 35771 26917
rect 35713 26908 35725 26911
rect 34848 26880 35725 26908
rect 34848 26868 34854 26880
rect 35713 26877 35725 26880
rect 35759 26877 35771 26911
rect 35713 26871 35771 26877
rect 34606 26840 34612 26852
rect 34532 26812 34612 26840
rect 34606 26800 34612 26812
rect 34664 26800 34670 26852
rect 34698 26800 34704 26852
rect 34756 26840 34762 26852
rect 36541 26843 36599 26849
rect 36541 26840 36553 26843
rect 34756 26812 36553 26840
rect 34756 26800 34762 26812
rect 36541 26809 36553 26812
rect 36587 26809 36599 26843
rect 36541 26803 36599 26809
rect 34790 26772 34796 26784
rect 34440 26744 34796 26772
rect 34790 26732 34796 26744
rect 34848 26732 34854 26784
rect 34977 26775 35035 26781
rect 34977 26741 34989 26775
rect 35023 26772 35035 26775
rect 35434 26772 35440 26784
rect 35023 26744 35440 26772
rect 35023 26741 35035 26744
rect 34977 26735 35035 26741
rect 35434 26732 35440 26744
rect 35492 26732 35498 26784
rect 35529 26775 35587 26781
rect 35529 26741 35541 26775
rect 35575 26772 35587 26775
rect 35618 26772 35624 26784
rect 35575 26744 35624 26772
rect 35575 26741 35587 26744
rect 35529 26735 35587 26741
rect 35618 26732 35624 26744
rect 35676 26732 35682 26784
rect 1104 26682 37628 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 37628 26682
rect 1104 26608 37628 26630
rect 7742 26568 7748 26580
rect 7703 26540 7748 26568
rect 7742 26528 7748 26540
rect 7800 26528 7806 26580
rect 8386 26528 8392 26580
rect 8444 26568 8450 26580
rect 8481 26571 8539 26577
rect 8481 26568 8493 26571
rect 8444 26540 8493 26568
rect 8444 26528 8450 26540
rect 8481 26537 8493 26540
rect 8527 26537 8539 26571
rect 8481 26531 8539 26537
rect 16301 26571 16359 26577
rect 16301 26537 16313 26571
rect 16347 26568 16359 26571
rect 18322 26568 18328 26580
rect 16347 26540 18328 26568
rect 16347 26537 16359 26540
rect 16301 26531 16359 26537
rect 18322 26528 18328 26540
rect 18380 26528 18386 26580
rect 18874 26568 18880 26580
rect 18835 26540 18880 26568
rect 18874 26528 18880 26540
rect 18932 26528 18938 26580
rect 18966 26528 18972 26580
rect 19024 26568 19030 26580
rect 22370 26568 22376 26580
rect 19024 26540 22376 26568
rect 19024 26528 19030 26540
rect 22370 26528 22376 26540
rect 22428 26528 22434 26580
rect 22465 26571 22523 26577
rect 22465 26537 22477 26571
rect 22511 26568 22523 26571
rect 22646 26568 22652 26580
rect 22511 26540 22652 26568
rect 22511 26537 22523 26540
rect 22465 26531 22523 26537
rect 22646 26528 22652 26540
rect 22704 26528 22710 26580
rect 24946 26528 24952 26580
rect 25004 26568 25010 26580
rect 25004 26540 26832 26568
rect 25004 26528 25010 26540
rect 10042 26460 10048 26512
rect 10100 26500 10106 26512
rect 10502 26500 10508 26512
rect 10100 26472 10508 26500
rect 10100 26460 10106 26472
rect 10502 26460 10508 26472
rect 10560 26460 10566 26512
rect 11333 26503 11391 26509
rect 11333 26469 11345 26503
rect 11379 26500 11391 26503
rect 16761 26503 16819 26509
rect 11379 26472 11928 26500
rect 11379 26469 11391 26472
rect 11333 26463 11391 26469
rect 10321 26435 10379 26441
rect 10321 26401 10333 26435
rect 10367 26401 10379 26435
rect 10321 26395 10379 26401
rect 7926 26364 7932 26376
rect 7887 26336 7932 26364
rect 7926 26324 7932 26336
rect 7984 26324 7990 26376
rect 8389 26367 8447 26373
rect 8389 26333 8401 26367
rect 8435 26364 8447 26367
rect 8754 26364 8760 26376
rect 8435 26336 8760 26364
rect 8435 26333 8447 26336
rect 8389 26327 8447 26333
rect 8754 26324 8760 26336
rect 8812 26324 8818 26376
rect 10042 26364 10048 26376
rect 10003 26336 10048 26364
rect 10042 26324 10048 26336
rect 10100 26324 10106 26376
rect 10336 26296 10364 26395
rect 11238 26392 11244 26444
rect 11296 26432 11302 26444
rect 11790 26432 11796 26444
rect 11296 26404 11796 26432
rect 11296 26392 11302 26404
rect 11790 26392 11796 26404
rect 11848 26392 11854 26444
rect 11900 26432 11928 26472
rect 16761 26469 16773 26503
rect 16807 26469 16819 26503
rect 19794 26500 19800 26512
rect 16761 26463 16819 26469
rect 17236 26472 19800 26500
rect 12069 26435 12127 26441
rect 12069 26432 12081 26435
rect 11900 26404 12081 26432
rect 12069 26401 12081 26404
rect 12115 26401 12127 26435
rect 12069 26395 12127 26401
rect 13078 26392 13084 26444
rect 13136 26432 13142 26444
rect 13541 26435 13599 26441
rect 13541 26432 13553 26435
rect 13136 26404 13553 26432
rect 13136 26392 13142 26404
rect 13541 26401 13553 26404
rect 13587 26432 13599 26435
rect 14921 26435 14979 26441
rect 14921 26432 14933 26435
rect 13587 26404 14933 26432
rect 13587 26401 13599 26404
rect 13541 26395 13599 26401
rect 14921 26401 14933 26404
rect 14967 26401 14979 26435
rect 15102 26432 15108 26444
rect 15063 26404 15108 26432
rect 14921 26395 14979 26401
rect 15102 26392 15108 26404
rect 15160 26392 15166 26444
rect 11146 26364 11152 26376
rect 11107 26336 11152 26364
rect 11146 26324 11152 26336
rect 11204 26324 11210 26376
rect 16117 26367 16175 26373
rect 16117 26333 16129 26367
rect 16163 26364 16175 26367
rect 16776 26364 16804 26463
rect 17236 26432 17264 26472
rect 19794 26460 19800 26472
rect 19852 26460 19858 26512
rect 19886 26460 19892 26512
rect 19944 26500 19950 26512
rect 23658 26500 23664 26512
rect 19944 26472 20116 26500
rect 19944 26460 19950 26472
rect 17402 26432 17408 26444
rect 17144 26404 17264 26432
rect 17315 26404 17408 26432
rect 17144 26373 17172 26404
rect 17402 26392 17408 26404
rect 17460 26432 17466 26444
rect 17460 26404 18184 26432
rect 17460 26392 17466 26404
rect 16163 26336 16804 26364
rect 17129 26367 17187 26373
rect 16163 26333 16175 26336
rect 16117 26327 16175 26333
rect 17129 26333 17141 26367
rect 17175 26333 17187 26367
rect 17129 26327 17187 26333
rect 17221 26367 17279 26373
rect 17221 26333 17233 26367
rect 17267 26364 17279 26367
rect 17586 26364 17592 26376
rect 17267 26336 17592 26364
rect 17267 26333 17279 26336
rect 17221 26327 17279 26333
rect 17586 26324 17592 26336
rect 17644 26324 17650 26376
rect 18156 26364 18184 26404
rect 18230 26392 18236 26444
rect 18288 26432 18294 26444
rect 18288 26404 18333 26432
rect 18288 26392 18294 26404
rect 18414 26392 18420 26444
rect 18472 26432 18478 26444
rect 20088 26441 20116 26472
rect 22066 26472 23664 26500
rect 19981 26435 20039 26441
rect 19981 26432 19993 26435
rect 18472 26404 19993 26432
rect 18472 26392 18478 26404
rect 19981 26401 19993 26404
rect 20027 26401 20039 26435
rect 19981 26395 20039 26401
rect 20073 26435 20131 26441
rect 20073 26401 20085 26435
rect 20119 26401 20131 26435
rect 20073 26395 20131 26401
rect 20622 26392 20628 26444
rect 20680 26392 20686 26444
rect 20717 26435 20775 26441
rect 20717 26401 20729 26435
rect 20763 26432 20775 26435
rect 22066 26432 22094 26472
rect 23658 26460 23664 26472
rect 23716 26460 23722 26512
rect 23937 26503 23995 26509
rect 23937 26469 23949 26503
rect 23983 26469 23995 26503
rect 23937 26463 23995 26469
rect 26605 26503 26663 26509
rect 26605 26469 26617 26503
rect 26651 26469 26663 26503
rect 26804 26500 26832 26540
rect 26878 26528 26884 26580
rect 26936 26568 26942 26580
rect 27157 26571 27215 26577
rect 27157 26568 27169 26571
rect 26936 26540 27169 26568
rect 26936 26528 26942 26540
rect 27157 26537 27169 26540
rect 27203 26537 27215 26571
rect 27157 26531 27215 26537
rect 28442 26528 28448 26580
rect 28500 26568 28506 26580
rect 28721 26571 28779 26577
rect 28721 26568 28733 26571
rect 28500 26540 28733 26568
rect 28500 26528 28506 26540
rect 28721 26537 28733 26540
rect 28767 26568 28779 26571
rect 30193 26571 30251 26577
rect 30193 26568 30205 26571
rect 28767 26540 30205 26568
rect 28767 26537 28779 26540
rect 28721 26531 28779 26537
rect 30193 26537 30205 26540
rect 30239 26568 30251 26571
rect 30466 26568 30472 26580
rect 30239 26540 30472 26568
rect 30239 26537 30251 26540
rect 30193 26531 30251 26537
rect 30466 26528 30472 26540
rect 30524 26528 30530 26580
rect 32306 26568 32312 26580
rect 30668 26540 32312 26568
rect 30668 26512 30696 26540
rect 32306 26528 32312 26540
rect 32364 26528 32370 26580
rect 34238 26568 34244 26580
rect 34199 26540 34244 26568
rect 34238 26528 34244 26540
rect 34296 26528 34302 26580
rect 35802 26528 35808 26580
rect 35860 26568 35866 26580
rect 37047 26571 37105 26577
rect 37047 26568 37059 26571
rect 35860 26540 37059 26568
rect 35860 26528 35866 26540
rect 37047 26537 37059 26540
rect 37093 26537 37105 26571
rect 37047 26531 37105 26537
rect 30650 26500 30656 26512
rect 26804 26472 30656 26500
rect 26605 26463 26663 26469
rect 20763 26404 22094 26432
rect 23385 26435 23443 26441
rect 20763 26401 20775 26404
rect 20717 26395 20775 26401
rect 23385 26401 23397 26435
rect 23431 26432 23443 26435
rect 23474 26432 23480 26444
rect 23431 26404 23480 26432
rect 23431 26401 23443 26404
rect 23385 26395 23443 26401
rect 23474 26392 23480 26404
rect 23532 26432 23538 26444
rect 23750 26432 23756 26444
rect 23532 26404 23756 26432
rect 23532 26392 23538 26404
rect 23750 26392 23756 26404
rect 23808 26392 23814 26444
rect 20640 26364 20668 26392
rect 18156 26336 20668 26364
rect 22094 26324 22100 26376
rect 22152 26324 22158 26376
rect 23569 26367 23627 26373
rect 23569 26333 23581 26367
rect 23615 26364 23627 26367
rect 23842 26364 23848 26376
rect 23615 26336 23848 26364
rect 23615 26333 23627 26336
rect 23569 26327 23627 26333
rect 23842 26324 23848 26336
rect 23900 26324 23906 26376
rect 23952 26364 23980 26463
rect 24670 26392 24676 26444
rect 24728 26432 24734 26444
rect 26053 26435 26111 26441
rect 24728 26404 25452 26432
rect 24728 26392 24734 26404
rect 25424 26373 25452 26404
rect 26053 26401 26065 26435
rect 26099 26432 26111 26435
rect 26234 26432 26240 26444
rect 26099 26404 26240 26432
rect 26099 26401 26111 26404
rect 26053 26395 26111 26401
rect 26234 26392 26240 26404
rect 26292 26392 26298 26444
rect 26620 26432 26648 26463
rect 30650 26460 30656 26472
rect 30708 26460 30714 26512
rect 33410 26500 33416 26512
rect 32692 26472 33416 26500
rect 31662 26432 31668 26444
rect 26620 26404 27936 26432
rect 31623 26404 31668 26432
rect 24765 26367 24823 26373
rect 24765 26364 24777 26367
rect 23952 26336 24777 26364
rect 24765 26333 24777 26336
rect 24811 26333 24823 26367
rect 24765 26327 24823 26333
rect 25409 26367 25467 26373
rect 25409 26333 25421 26367
rect 25455 26333 25467 26367
rect 25409 26327 25467 26333
rect 27249 26367 27307 26373
rect 27249 26333 27261 26367
rect 27295 26364 27307 26367
rect 27338 26364 27344 26376
rect 27295 26336 27344 26364
rect 27295 26333 27307 26336
rect 27249 26327 27307 26333
rect 27338 26324 27344 26336
rect 27396 26324 27402 26376
rect 27908 26373 27936 26404
rect 31662 26392 31668 26404
rect 31720 26392 31726 26444
rect 32692 26441 32720 26472
rect 33410 26460 33416 26472
rect 33468 26460 33474 26512
rect 34606 26500 34612 26512
rect 34440 26472 34612 26500
rect 32677 26435 32735 26441
rect 32677 26401 32689 26435
rect 32723 26401 32735 26435
rect 32677 26395 32735 26401
rect 27893 26367 27951 26373
rect 27893 26333 27905 26367
rect 27939 26333 27951 26367
rect 28626 26364 28632 26376
rect 27893 26327 27951 26333
rect 28368 26336 28632 26364
rect 11330 26296 11336 26308
rect 10336 26268 11336 26296
rect 11330 26256 11336 26268
rect 11388 26256 11394 26308
rect 11422 26256 11428 26308
rect 11480 26296 11486 26308
rect 14829 26299 14887 26305
rect 11480 26268 12558 26296
rect 11480 26256 11486 26268
rect 14829 26265 14841 26299
rect 14875 26296 14887 26299
rect 20990 26296 20996 26308
rect 14875 26268 20852 26296
rect 20951 26268 20996 26296
rect 14875 26265 14887 26268
rect 14829 26259 14887 26265
rect 9674 26228 9680 26240
rect 9635 26200 9680 26228
rect 9674 26188 9680 26200
rect 9732 26188 9738 26240
rect 10134 26228 10140 26240
rect 10095 26200 10140 26228
rect 10134 26188 10140 26200
rect 10192 26188 10198 26240
rect 13814 26188 13820 26240
rect 13872 26228 13878 26240
rect 14461 26231 14519 26237
rect 14461 26228 14473 26231
rect 13872 26200 14473 26228
rect 13872 26188 13878 26200
rect 14461 26197 14473 26200
rect 14507 26197 14519 26231
rect 14461 26191 14519 26197
rect 18506 26188 18512 26240
rect 18564 26228 18570 26240
rect 19518 26228 19524 26240
rect 18564 26200 18609 26228
rect 19479 26200 19524 26228
rect 18564 26188 18570 26200
rect 19518 26188 19524 26200
rect 19576 26188 19582 26240
rect 19886 26228 19892 26240
rect 19847 26200 19892 26228
rect 19886 26188 19892 26200
rect 19944 26188 19950 26240
rect 20824 26228 20852 26268
rect 20990 26256 20996 26268
rect 21048 26256 21054 26308
rect 25314 26296 25320 26308
rect 22296 26268 25176 26296
rect 25275 26268 25320 26296
rect 22296 26228 22324 26268
rect 23474 26228 23480 26240
rect 20824 26200 22324 26228
rect 23435 26200 23480 26228
rect 23474 26188 23480 26200
rect 23532 26188 23538 26240
rect 24578 26228 24584 26240
rect 24539 26200 24584 26228
rect 24578 26188 24584 26200
rect 24636 26188 24642 26240
rect 25148 26228 25176 26268
rect 25314 26256 25320 26268
rect 25372 26256 25378 26308
rect 28368 26296 28396 26336
rect 28626 26324 28632 26336
rect 28684 26324 28690 26376
rect 31938 26324 31944 26376
rect 31996 26364 32002 26376
rect 32692 26364 32720 26395
rect 33042 26392 33048 26444
rect 33100 26392 33106 26444
rect 33870 26432 33876 26444
rect 33831 26404 33876 26432
rect 33870 26392 33876 26404
rect 33928 26392 33934 26444
rect 32950 26364 32956 26376
rect 31996 26336 32041 26364
rect 32140 26336 32720 26364
rect 32911 26336 32956 26364
rect 31996 26324 32002 26336
rect 28534 26296 28540 26308
rect 25424 26268 28396 26296
rect 28495 26268 28540 26296
rect 25424 26228 25452 26268
rect 28534 26256 28540 26268
rect 28592 26256 28598 26308
rect 28644 26296 28672 26324
rect 28737 26299 28795 26305
rect 28737 26296 28749 26299
rect 28644 26268 28749 26296
rect 28737 26265 28749 26268
rect 28783 26265 28795 26299
rect 28737 26259 28795 26265
rect 31202 26256 31208 26308
rect 31260 26256 31266 26308
rect 32140 26296 32168 26336
rect 32950 26324 32956 26336
rect 33008 26324 33014 26376
rect 31956 26268 32168 26296
rect 25148 26200 25452 26228
rect 26050 26188 26056 26240
rect 26108 26228 26114 26240
rect 26145 26231 26203 26237
rect 26145 26228 26157 26231
rect 26108 26200 26157 26228
rect 26108 26188 26114 26200
rect 26145 26197 26157 26200
rect 26191 26197 26203 26231
rect 26145 26191 26203 26197
rect 26237 26231 26295 26237
rect 26237 26197 26249 26231
rect 26283 26228 26295 26231
rect 26326 26228 26332 26240
rect 26283 26200 26332 26228
rect 26283 26197 26295 26200
rect 26237 26191 26295 26197
rect 26326 26188 26332 26200
rect 26384 26188 26390 26240
rect 27706 26228 27712 26240
rect 27667 26200 27712 26228
rect 27706 26188 27712 26200
rect 27764 26188 27770 26240
rect 28902 26228 28908 26240
rect 28863 26200 28908 26228
rect 28902 26188 28908 26200
rect 28960 26188 28966 26240
rect 31294 26188 31300 26240
rect 31352 26228 31358 26240
rect 31956 26228 31984 26268
rect 32582 26256 32588 26308
rect 32640 26296 32646 26308
rect 33060 26305 33088 26392
rect 33134 26324 33140 26376
rect 33192 26364 33198 26376
rect 33962 26364 33968 26376
rect 33192 26336 33237 26364
rect 33923 26336 33968 26364
rect 33192 26324 33198 26336
rect 33962 26324 33968 26336
rect 34020 26324 34026 26376
rect 34440 26364 34468 26472
rect 34606 26460 34612 26472
rect 34664 26460 34670 26512
rect 34514 26392 34520 26444
rect 34572 26432 34578 26444
rect 35253 26435 35311 26441
rect 35253 26432 35265 26435
rect 34572 26404 35265 26432
rect 34572 26392 34578 26404
rect 35253 26401 35265 26404
rect 35299 26432 35311 26435
rect 35618 26432 35624 26444
rect 35299 26404 35388 26432
rect 35579 26404 35624 26432
rect 35299 26401 35311 26404
rect 35253 26395 35311 26401
rect 35360 26376 35388 26404
rect 35618 26392 35624 26404
rect 35676 26392 35682 26444
rect 34440 26336 34560 26364
rect 34532 26308 34560 26336
rect 35342 26324 35348 26376
rect 35400 26324 35406 26376
rect 32815 26299 32873 26305
rect 32815 26296 32827 26299
rect 32640 26268 32827 26296
rect 32640 26256 32646 26268
rect 32815 26265 32827 26268
rect 32861 26265 32873 26299
rect 32815 26259 32873 26265
rect 33045 26299 33103 26305
rect 33045 26265 33057 26299
rect 33091 26265 33103 26299
rect 33045 26259 33103 26265
rect 34514 26256 34520 26308
rect 34572 26256 34578 26308
rect 36446 26256 36452 26308
rect 36504 26256 36510 26308
rect 31352 26200 31984 26228
rect 33321 26231 33379 26237
rect 31352 26188 31358 26200
rect 33321 26197 33333 26231
rect 33367 26228 33379 26231
rect 33686 26228 33692 26240
rect 33367 26200 33692 26228
rect 33367 26197 33379 26200
rect 33321 26191 33379 26197
rect 33686 26188 33692 26200
rect 33744 26188 33750 26240
rect 1104 26138 37628 26160
rect 1104 26086 4874 26138
rect 4926 26086 4938 26138
rect 4990 26086 5002 26138
rect 5054 26086 5066 26138
rect 5118 26086 5130 26138
rect 5182 26086 35594 26138
rect 35646 26086 35658 26138
rect 35710 26086 35722 26138
rect 35774 26086 35786 26138
rect 35838 26086 35850 26138
rect 35902 26086 37628 26138
rect 1104 26064 37628 26086
rect 9048 25996 10916 26024
rect 8389 25891 8447 25897
rect 8389 25857 8401 25891
rect 8435 25888 8447 25891
rect 9048 25888 9076 25996
rect 9766 25956 9772 25968
rect 9232 25928 9772 25956
rect 8435 25860 9076 25888
rect 8435 25857 8447 25860
rect 8389 25851 8447 25857
rect 9122 25848 9128 25900
rect 9180 25888 9186 25900
rect 9232 25897 9260 25928
rect 9766 25916 9772 25928
rect 9824 25916 9830 25968
rect 9950 25916 9956 25968
rect 10008 25916 10014 25968
rect 10888 25900 10916 25996
rect 12802 25984 12808 26036
rect 12860 26024 12866 26036
rect 15657 26027 15715 26033
rect 15657 26024 15669 26027
rect 12860 25996 15669 26024
rect 12860 25984 12866 25996
rect 15657 25993 15669 25996
rect 15703 25993 15715 26027
rect 15657 25987 15715 25993
rect 19245 26027 19303 26033
rect 19245 25993 19257 26027
rect 19291 25993 19303 26027
rect 19245 25987 19303 25993
rect 14182 25956 14188 25968
rect 14143 25928 14188 25956
rect 14182 25916 14188 25928
rect 14240 25916 14246 25968
rect 15194 25916 15200 25968
rect 15252 25916 15258 25968
rect 18322 25956 18328 25968
rect 18283 25928 18328 25956
rect 18322 25916 18328 25928
rect 18380 25916 18386 25968
rect 19260 25956 19288 25987
rect 19702 25984 19708 26036
rect 19760 26024 19766 26036
rect 19760 25996 22140 26024
rect 19760 25984 19766 25996
rect 19981 25959 20039 25965
rect 19981 25956 19993 25959
rect 19260 25928 19993 25956
rect 19981 25925 19993 25928
rect 20027 25925 20039 25959
rect 19981 25919 20039 25925
rect 20990 25916 20996 25968
rect 21048 25916 21054 25968
rect 9217 25891 9275 25897
rect 9217 25888 9229 25891
rect 9180 25860 9229 25888
rect 9180 25848 9186 25860
rect 9217 25857 9229 25860
rect 9263 25857 9275 25891
rect 9217 25851 9275 25857
rect 10870 25848 10876 25900
rect 10928 25888 10934 25900
rect 12161 25891 12219 25897
rect 12161 25888 12173 25891
rect 10928 25860 12173 25888
rect 10928 25848 10934 25860
rect 12161 25857 12173 25860
rect 12207 25857 12219 25891
rect 12161 25851 12219 25857
rect 13265 25891 13323 25897
rect 13265 25857 13277 25891
rect 13311 25888 13323 25891
rect 13814 25888 13820 25900
rect 13311 25860 13820 25888
rect 13311 25857 13323 25860
rect 13265 25851 13323 25857
rect 13814 25848 13820 25860
rect 13872 25848 13878 25900
rect 16117 25891 16175 25897
rect 16117 25857 16129 25891
rect 16163 25857 16175 25891
rect 16117 25851 16175 25857
rect 8570 25780 8576 25832
rect 8628 25820 8634 25832
rect 9493 25823 9551 25829
rect 9493 25820 9505 25823
rect 8628 25792 9505 25820
rect 8628 25780 8634 25792
rect 9493 25789 9505 25792
rect 9539 25789 9551 25823
rect 9493 25783 9551 25789
rect 13722 25780 13728 25832
rect 13780 25820 13786 25832
rect 13909 25823 13967 25829
rect 13909 25820 13921 25823
rect 13780 25792 13921 25820
rect 13780 25780 13786 25792
rect 13909 25789 13921 25792
rect 13955 25789 13967 25823
rect 15654 25820 15660 25832
rect 13909 25783 13967 25789
rect 14016 25792 15660 25820
rect 10502 25712 10508 25764
rect 10560 25752 10566 25764
rect 10965 25755 11023 25761
rect 10965 25752 10977 25755
rect 10560 25724 10977 25752
rect 10560 25712 10566 25724
rect 10965 25721 10977 25724
rect 11011 25752 11023 25755
rect 14016 25752 14044 25792
rect 15654 25780 15660 25792
rect 15712 25780 15718 25832
rect 16132 25820 16160 25851
rect 17218 25848 17224 25900
rect 17276 25848 17282 25900
rect 19061 25891 19119 25897
rect 19061 25857 19073 25891
rect 19107 25888 19119 25891
rect 19518 25888 19524 25900
rect 19107 25860 19524 25888
rect 19107 25857 19119 25860
rect 19061 25851 19119 25857
rect 19518 25848 19524 25860
rect 19576 25848 19582 25900
rect 22112 25897 22140 25996
rect 23750 25984 23756 26036
rect 23808 26024 23814 26036
rect 26050 26024 26056 26036
rect 23808 25996 26056 26024
rect 23808 25984 23814 25996
rect 26050 25984 26056 25996
rect 26108 25984 26114 26036
rect 26145 26027 26203 26033
rect 26145 25993 26157 26027
rect 26191 26024 26203 26027
rect 28350 26024 28356 26036
rect 26191 25996 28356 26024
rect 26191 25993 26203 25996
rect 26145 25987 26203 25993
rect 28350 25984 28356 25996
rect 28408 25984 28414 26036
rect 30469 26027 30527 26033
rect 30469 25993 30481 26027
rect 30515 25993 30527 26027
rect 32030 26024 32036 26036
rect 30469 25987 30527 25993
rect 30576 25996 32036 26024
rect 25314 25956 25320 25968
rect 23598 25928 25320 25956
rect 25314 25916 25320 25928
rect 25372 25916 25378 25968
rect 26326 25956 26332 25968
rect 25516 25928 26332 25956
rect 22097 25891 22155 25897
rect 22097 25857 22109 25891
rect 22143 25857 22155 25891
rect 22097 25851 22155 25857
rect 24762 25848 24768 25900
rect 24820 25888 24826 25900
rect 24857 25891 24915 25897
rect 24857 25888 24869 25891
rect 24820 25860 24869 25888
rect 24820 25848 24826 25860
rect 24857 25857 24869 25860
rect 24903 25857 24915 25891
rect 24857 25851 24915 25857
rect 24949 25891 25007 25897
rect 24949 25857 24961 25891
rect 24995 25888 25007 25891
rect 25516 25888 25544 25928
rect 26326 25916 26332 25928
rect 26384 25916 26390 25968
rect 27433 25959 27491 25965
rect 27433 25925 27445 25959
rect 27479 25956 27491 25959
rect 27706 25956 27712 25968
rect 27479 25928 27712 25956
rect 27479 25925 27491 25928
rect 27433 25919 27491 25925
rect 27706 25916 27712 25928
rect 27764 25916 27770 25968
rect 27890 25916 27896 25968
rect 27948 25916 27954 25968
rect 30484 25956 30512 25987
rect 30576 25965 30604 25996
rect 32030 25984 32036 25996
rect 32088 25984 32094 26036
rect 33505 26027 33563 26033
rect 33505 25993 33517 26027
rect 33551 26024 33563 26027
rect 33870 26024 33876 26036
rect 33551 25996 33876 26024
rect 33551 25993 33563 25996
rect 33505 25987 33563 25993
rect 33870 25984 33876 25996
rect 33928 25984 33934 26036
rect 29840 25928 30512 25956
rect 30561 25959 30619 25965
rect 24995 25860 25544 25888
rect 25608 25860 26280 25888
rect 24995 25857 25007 25860
rect 24949 25851 25007 25857
rect 16132 25792 18552 25820
rect 11011 25724 14044 25752
rect 18524 25752 18552 25792
rect 18598 25780 18604 25832
rect 18656 25820 18662 25832
rect 19702 25820 19708 25832
rect 18656 25792 18701 25820
rect 19663 25792 19708 25820
rect 18656 25780 18662 25792
rect 19702 25780 19708 25792
rect 19760 25780 19766 25832
rect 22373 25823 22431 25829
rect 22373 25789 22385 25823
rect 22419 25820 22431 25823
rect 24578 25820 24584 25832
rect 22419 25792 24584 25820
rect 22419 25789 22431 25792
rect 22373 25783 22431 25789
rect 24578 25780 24584 25792
rect 24636 25780 24642 25832
rect 19426 25752 19432 25764
rect 18524 25724 19432 25752
rect 11011 25721 11023 25724
rect 10965 25715 11023 25721
rect 19426 25712 19432 25724
rect 19484 25712 19490 25764
rect 23474 25712 23480 25764
rect 23532 25752 23538 25764
rect 23845 25755 23903 25761
rect 23845 25752 23857 25755
rect 23532 25724 23857 25752
rect 23532 25712 23538 25724
rect 23845 25721 23857 25724
rect 23891 25752 23903 25755
rect 24780 25752 24808 25848
rect 25608 25832 25636 25860
rect 25133 25823 25191 25829
rect 25133 25789 25145 25823
rect 25179 25820 25191 25823
rect 25590 25820 25596 25832
rect 25179 25792 25596 25820
rect 25179 25789 25191 25792
rect 25133 25783 25191 25789
rect 25590 25780 25596 25792
rect 25648 25780 25654 25832
rect 26252 25829 26280 25860
rect 26237 25823 26295 25829
rect 26237 25789 26249 25823
rect 26283 25789 26295 25823
rect 26237 25783 26295 25789
rect 23891 25724 24808 25752
rect 23891 25721 23903 25724
rect 23845 25715 23903 25721
rect 8478 25684 8484 25696
rect 8439 25656 8484 25684
rect 8478 25644 8484 25656
rect 8536 25644 8542 25696
rect 12158 25644 12164 25696
rect 12216 25684 12222 25696
rect 12253 25687 12311 25693
rect 12253 25684 12265 25687
rect 12216 25656 12265 25684
rect 12216 25644 12222 25656
rect 12253 25653 12265 25656
rect 12299 25653 12311 25687
rect 12253 25647 12311 25653
rect 13449 25687 13507 25693
rect 13449 25653 13461 25687
rect 13495 25684 13507 25687
rect 14550 25684 14556 25696
rect 13495 25656 14556 25684
rect 13495 25653 13507 25656
rect 13449 25647 13507 25653
rect 14550 25644 14556 25656
rect 14608 25644 14614 25696
rect 16298 25684 16304 25696
rect 16259 25656 16304 25684
rect 16298 25644 16304 25656
rect 16356 25644 16362 25696
rect 16574 25644 16580 25696
rect 16632 25684 16638 25696
rect 16853 25687 16911 25693
rect 16853 25684 16865 25687
rect 16632 25656 16865 25684
rect 16632 25644 16638 25656
rect 16853 25653 16865 25656
rect 16899 25653 16911 25687
rect 16853 25647 16911 25653
rect 19978 25644 19984 25696
rect 20036 25684 20042 25696
rect 21082 25684 21088 25696
rect 20036 25656 21088 25684
rect 20036 25644 20042 25656
rect 21082 25644 21088 25656
rect 21140 25684 21146 25696
rect 21453 25687 21511 25693
rect 21453 25684 21465 25687
rect 21140 25656 21465 25684
rect 21140 25644 21146 25656
rect 21453 25653 21465 25656
rect 21499 25653 21511 25687
rect 24486 25684 24492 25696
rect 24447 25656 24492 25684
rect 21453 25647 21511 25653
rect 24486 25644 24492 25656
rect 24544 25644 24550 25696
rect 24946 25644 24952 25696
rect 25004 25684 25010 25696
rect 25685 25687 25743 25693
rect 25685 25684 25697 25687
rect 25004 25656 25697 25684
rect 25004 25644 25010 25656
rect 25685 25653 25697 25656
rect 25731 25653 25743 25687
rect 26344 25684 26372 25916
rect 29549 25891 29607 25897
rect 29549 25857 29561 25891
rect 29595 25857 29607 25891
rect 29549 25851 29607 25857
rect 29641 25891 29699 25897
rect 29641 25857 29653 25891
rect 29687 25888 29699 25891
rect 29730 25888 29736 25900
rect 29687 25860 29736 25888
rect 29687 25857 29699 25860
rect 29641 25851 29699 25857
rect 27154 25820 27160 25832
rect 27115 25792 27160 25820
rect 27154 25780 27160 25792
rect 27212 25780 27218 25832
rect 29564 25820 29592 25851
rect 29730 25848 29736 25860
rect 29788 25848 29794 25900
rect 29840 25897 29868 25928
rect 30561 25925 30573 25959
rect 30607 25925 30619 25959
rect 30561 25919 30619 25925
rect 29825 25891 29883 25897
rect 29825 25857 29837 25891
rect 29871 25857 29883 25891
rect 29825 25851 29883 25857
rect 30377 25891 30435 25897
rect 30377 25857 30389 25891
rect 30423 25888 30435 25891
rect 30466 25888 30472 25900
rect 30423 25860 30472 25888
rect 30423 25857 30435 25860
rect 30377 25851 30435 25857
rect 30466 25848 30472 25860
rect 30524 25848 30530 25900
rect 30576 25820 30604 25919
rect 31570 25916 31576 25968
rect 31628 25956 31634 25968
rect 31628 25928 32536 25956
rect 31628 25916 31634 25928
rect 30650 25848 30656 25900
rect 30708 25888 30714 25900
rect 31110 25888 31116 25900
rect 30708 25860 30753 25888
rect 31071 25860 31116 25888
rect 30708 25848 30714 25860
rect 31110 25848 31116 25860
rect 31168 25848 31174 25900
rect 31294 25888 31300 25900
rect 31255 25860 31300 25888
rect 31294 25848 31300 25860
rect 31352 25848 31358 25900
rect 32508 25897 32536 25928
rect 33042 25916 33048 25968
rect 33100 25956 33106 25968
rect 33413 25959 33471 25965
rect 33413 25956 33425 25959
rect 33100 25928 33425 25956
rect 33100 25916 33106 25928
rect 33413 25925 33425 25928
rect 33459 25925 33471 25959
rect 36262 25956 36268 25968
rect 35742 25928 36268 25956
rect 33413 25919 33471 25925
rect 36262 25916 36268 25928
rect 36320 25916 36326 25968
rect 32493 25891 32551 25897
rect 32493 25857 32505 25891
rect 32539 25857 32551 25891
rect 32493 25851 32551 25857
rect 32582 25848 32588 25900
rect 32640 25888 32646 25900
rect 32769 25891 32827 25897
rect 32640 25860 32685 25888
rect 32640 25848 32646 25860
rect 32769 25857 32781 25891
rect 32815 25857 32827 25891
rect 32769 25851 32827 25857
rect 29564 25792 30604 25820
rect 31754 25780 31760 25832
rect 31812 25820 31818 25832
rect 32784 25820 32812 25851
rect 33134 25848 33140 25900
rect 33192 25888 33198 25900
rect 33318 25888 33324 25900
rect 33192 25860 33324 25888
rect 33192 25848 33198 25860
rect 33318 25848 33324 25860
rect 33376 25848 33382 25900
rect 33781 25891 33839 25897
rect 33781 25857 33793 25891
rect 33827 25888 33839 25891
rect 34606 25888 34612 25900
rect 33827 25860 34612 25888
rect 33827 25857 33839 25860
rect 33781 25851 33839 25857
rect 34606 25848 34612 25860
rect 34664 25848 34670 25900
rect 36170 25820 36176 25832
rect 31812 25792 32812 25820
rect 36131 25792 36176 25820
rect 31812 25780 31818 25792
rect 36170 25780 36176 25792
rect 36228 25780 36234 25832
rect 36449 25823 36507 25829
rect 36449 25789 36461 25823
rect 36495 25789 36507 25823
rect 36449 25783 36507 25789
rect 29733 25755 29791 25761
rect 29733 25721 29745 25755
rect 29779 25752 29791 25755
rect 32309 25755 32367 25761
rect 32309 25752 32321 25755
rect 29779 25724 32321 25752
rect 29779 25721 29791 25724
rect 29733 25715 29791 25721
rect 32309 25721 32321 25724
rect 32355 25721 32367 25755
rect 32309 25715 32367 25721
rect 32398 25712 32404 25764
rect 32456 25752 32462 25764
rect 34514 25752 34520 25764
rect 32456 25724 34520 25752
rect 32456 25712 32462 25724
rect 34514 25712 34520 25724
rect 34572 25752 34578 25764
rect 34701 25755 34759 25761
rect 34701 25752 34713 25755
rect 34572 25724 34713 25752
rect 34572 25712 34578 25724
rect 34701 25721 34713 25724
rect 34747 25721 34759 25755
rect 34701 25715 34759 25721
rect 28905 25687 28963 25693
rect 28905 25684 28917 25687
rect 26344 25656 28917 25684
rect 25685 25647 25743 25653
rect 28905 25653 28917 25656
rect 28951 25684 28963 25687
rect 28994 25684 29000 25696
rect 28951 25656 29000 25684
rect 28951 25653 28963 25656
rect 28905 25647 28963 25653
rect 28994 25644 29000 25656
rect 29052 25644 29058 25696
rect 29362 25684 29368 25696
rect 29323 25656 29368 25684
rect 29362 25644 29368 25656
rect 29420 25644 29426 25696
rect 30374 25644 30380 25696
rect 30432 25684 30438 25696
rect 31205 25687 31263 25693
rect 31205 25684 31217 25687
rect 30432 25656 31217 25684
rect 30432 25644 30438 25656
rect 31205 25653 31217 25656
rect 31251 25653 31263 25687
rect 32766 25684 32772 25696
rect 32727 25656 32772 25684
rect 31205 25647 31263 25653
rect 32766 25644 32772 25656
rect 32824 25644 32830 25696
rect 35434 25644 35440 25696
rect 35492 25684 35498 25696
rect 36464 25684 36492 25783
rect 35492 25656 36492 25684
rect 35492 25644 35498 25656
rect 1104 25594 37628 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 37628 25594
rect 1104 25520 37628 25542
rect 8570 25480 8576 25492
rect 8531 25452 8576 25480
rect 8570 25440 8576 25452
rect 8628 25440 8634 25492
rect 12066 25440 12072 25492
rect 12124 25480 12130 25492
rect 12897 25483 12955 25489
rect 12897 25480 12909 25483
rect 12124 25452 12909 25480
rect 12124 25440 12130 25452
rect 12897 25449 12909 25452
rect 12943 25480 12955 25483
rect 18325 25483 18383 25489
rect 18325 25480 18337 25483
rect 12943 25452 18337 25480
rect 12943 25449 12955 25452
rect 12897 25443 12955 25449
rect 18325 25449 18337 25452
rect 18371 25449 18383 25483
rect 18325 25443 18383 25449
rect 18506 25440 18512 25492
rect 18564 25480 18570 25492
rect 19429 25483 19487 25489
rect 19429 25480 19441 25483
rect 18564 25452 19441 25480
rect 18564 25440 18570 25452
rect 19429 25449 19441 25452
rect 19475 25449 19487 25483
rect 19429 25443 19487 25449
rect 20901 25483 20959 25489
rect 20901 25449 20913 25483
rect 20947 25480 20959 25483
rect 20990 25480 20996 25492
rect 20947 25452 20996 25480
rect 20947 25449 20959 25452
rect 20901 25443 20959 25449
rect 20990 25440 20996 25452
rect 21048 25440 21054 25492
rect 28350 25480 28356 25492
rect 28311 25452 28356 25480
rect 28350 25440 28356 25452
rect 28408 25440 28414 25492
rect 29730 25440 29736 25492
rect 29788 25480 29794 25492
rect 31110 25480 31116 25492
rect 29788 25452 31116 25480
rect 29788 25440 29794 25452
rect 31110 25440 31116 25452
rect 31168 25440 31174 25492
rect 31478 25480 31484 25492
rect 31439 25452 31484 25480
rect 31478 25440 31484 25452
rect 31536 25440 31542 25492
rect 31754 25480 31760 25492
rect 31715 25452 31760 25480
rect 31754 25440 31760 25452
rect 31812 25440 31818 25492
rect 32582 25480 32588 25492
rect 32543 25452 32588 25480
rect 32582 25440 32588 25452
rect 32640 25440 32646 25492
rect 35897 25483 35955 25489
rect 35897 25449 35909 25483
rect 35943 25480 35955 25483
rect 36170 25480 36176 25492
rect 35943 25452 36176 25480
rect 35943 25449 35955 25452
rect 35897 25443 35955 25449
rect 36170 25440 36176 25452
rect 36228 25440 36234 25492
rect 36262 25440 36268 25492
rect 36320 25480 36326 25492
rect 36449 25483 36507 25489
rect 36449 25480 36461 25483
rect 36320 25452 36461 25480
rect 36320 25440 36326 25452
rect 36449 25449 36461 25452
rect 36495 25449 36507 25483
rect 36449 25443 36507 25449
rect 19334 25372 19340 25424
rect 19392 25412 19398 25424
rect 19392 25384 20116 25412
rect 19392 25372 19398 25384
rect 9582 25304 9588 25356
rect 9640 25344 9646 25356
rect 9861 25347 9919 25353
rect 9861 25344 9873 25347
rect 9640 25316 9873 25344
rect 9640 25304 9646 25316
rect 9861 25313 9873 25316
rect 9907 25313 9919 25347
rect 11146 25344 11152 25356
rect 11107 25316 11152 25344
rect 9861 25307 9919 25313
rect 11146 25304 11152 25316
rect 11204 25304 11210 25356
rect 14550 25344 14556 25356
rect 14511 25316 14556 25344
rect 14550 25304 14556 25316
rect 14608 25304 14614 25356
rect 14642 25304 14648 25356
rect 14700 25344 14706 25356
rect 14700 25316 16252 25344
rect 14700 25304 14706 25316
rect 7926 25276 7932 25288
rect 7887 25248 7932 25276
rect 7926 25236 7932 25248
rect 7984 25236 7990 25288
rect 8389 25279 8447 25285
rect 8389 25245 8401 25279
rect 8435 25276 8447 25279
rect 9674 25276 9680 25288
rect 8435 25248 9680 25276
rect 8435 25245 8447 25248
rect 8389 25239 8447 25245
rect 9674 25236 9680 25248
rect 9732 25236 9738 25288
rect 10505 25279 10563 25285
rect 10505 25245 10517 25279
rect 10551 25276 10563 25279
rect 10962 25276 10968 25288
rect 10551 25248 10968 25276
rect 10551 25245 10563 25248
rect 10505 25239 10563 25245
rect 10962 25236 10968 25248
rect 11020 25236 11026 25288
rect 13722 25236 13728 25288
rect 13780 25276 13786 25288
rect 14277 25279 14335 25285
rect 14277 25276 14289 25279
rect 13780 25248 14289 25276
rect 13780 25236 13786 25248
rect 14277 25245 14289 25248
rect 14323 25245 14335 25279
rect 16224 25276 16252 25316
rect 16298 25304 16304 25356
rect 16356 25344 16362 25356
rect 16853 25347 16911 25353
rect 16853 25344 16865 25347
rect 16356 25316 16865 25344
rect 16356 25304 16362 25316
rect 16853 25313 16865 25316
rect 16899 25313 16911 25347
rect 19886 25344 19892 25356
rect 19847 25316 19892 25344
rect 16853 25307 16911 25313
rect 19886 25304 19892 25316
rect 19944 25304 19950 25356
rect 20088 25353 20116 25384
rect 20073 25347 20131 25353
rect 20073 25313 20085 25347
rect 20119 25344 20131 25347
rect 20162 25344 20168 25356
rect 20119 25316 20168 25344
rect 20119 25313 20131 25316
rect 20073 25307 20131 25313
rect 20162 25304 20168 25316
rect 20220 25304 20226 25356
rect 23750 25344 23756 25356
rect 23711 25316 23756 25344
rect 23750 25304 23756 25316
rect 23808 25304 23814 25356
rect 23842 25304 23848 25356
rect 23900 25344 23906 25356
rect 24673 25347 24731 25353
rect 24673 25344 24685 25347
rect 23900 25316 24685 25344
rect 23900 25304 23906 25316
rect 24673 25313 24685 25316
rect 24719 25313 24731 25347
rect 24673 25307 24731 25313
rect 26605 25347 26663 25353
rect 26605 25313 26617 25347
rect 26651 25344 26663 25347
rect 26970 25344 26976 25356
rect 26651 25316 26976 25344
rect 26651 25313 26663 25316
rect 26605 25307 26663 25313
rect 26970 25304 26976 25316
rect 27028 25304 27034 25356
rect 30558 25344 30564 25356
rect 30519 25316 30564 25344
rect 30558 25304 30564 25316
rect 30616 25304 30622 25356
rect 30650 25304 30656 25356
rect 30708 25344 30714 25356
rect 31481 25347 31539 25353
rect 31481 25344 31493 25347
rect 30708 25316 31493 25344
rect 30708 25304 30714 25316
rect 31481 25313 31493 25316
rect 31527 25313 31539 25347
rect 31481 25307 31539 25313
rect 33597 25347 33655 25353
rect 33597 25313 33609 25347
rect 33643 25344 33655 25347
rect 33643 25316 35112 25344
rect 33643 25313 33655 25316
rect 33597 25307 33655 25313
rect 16577 25279 16635 25285
rect 16577 25276 16589 25279
rect 16224 25248 16589 25276
rect 14277 25239 14335 25245
rect 16577 25245 16589 25248
rect 16623 25245 16635 25279
rect 16577 25239 16635 25245
rect 8202 25168 8208 25220
rect 8260 25208 8266 25220
rect 11425 25211 11483 25217
rect 8260 25180 9720 25208
rect 8260 25168 8266 25180
rect 7742 25140 7748 25152
rect 7703 25112 7748 25140
rect 7742 25100 7748 25112
rect 7800 25100 7806 25152
rect 9306 25140 9312 25152
rect 9267 25112 9312 25140
rect 9306 25100 9312 25112
rect 9364 25100 9370 25152
rect 9692 25149 9720 25180
rect 11425 25177 11437 25211
rect 11471 25177 11483 25211
rect 11425 25171 11483 25177
rect 9677 25143 9735 25149
rect 9677 25109 9689 25143
rect 9723 25109 9735 25143
rect 9677 25103 9735 25109
rect 9769 25143 9827 25149
rect 9769 25109 9781 25143
rect 9815 25140 9827 25143
rect 10502 25140 10508 25152
rect 9815 25112 10508 25140
rect 9815 25109 9827 25112
rect 9769 25103 9827 25109
rect 10502 25100 10508 25112
rect 10560 25100 10566 25152
rect 10689 25143 10747 25149
rect 10689 25109 10701 25143
rect 10735 25140 10747 25143
rect 11440 25140 11468 25171
rect 12158 25168 12164 25220
rect 12216 25168 12222 25220
rect 14292 25208 14320 25239
rect 14642 25208 14648 25220
rect 14292 25180 14648 25208
rect 14642 25168 14648 25180
rect 14700 25168 14706 25220
rect 15286 25168 15292 25220
rect 15344 25168 15350 25220
rect 16592 25208 16620 25239
rect 17954 25236 17960 25288
rect 18012 25236 18018 25288
rect 20714 25236 20720 25288
rect 20772 25276 20778 25288
rect 20993 25279 21051 25285
rect 20993 25276 21005 25279
rect 20772 25248 21005 25276
rect 20772 25236 20778 25248
rect 20993 25245 21005 25248
rect 21039 25245 21051 25279
rect 20993 25239 21051 25245
rect 22649 25279 22707 25285
rect 22649 25245 22661 25279
rect 22695 25276 22707 25279
rect 23661 25279 23719 25285
rect 22695 25248 23336 25276
rect 22695 25245 22707 25248
rect 22649 25239 22707 25245
rect 16942 25208 16948 25220
rect 16592 25180 16948 25208
rect 16942 25168 16948 25180
rect 17000 25168 17006 25220
rect 10735 25112 11468 25140
rect 10735 25109 10747 25112
rect 10689 25103 10747 25109
rect 14366 25100 14372 25152
rect 14424 25140 14430 25152
rect 15930 25140 15936 25152
rect 14424 25112 15936 25140
rect 14424 25100 14430 25112
rect 15930 25100 15936 25112
rect 15988 25140 15994 25152
rect 16025 25143 16083 25149
rect 16025 25140 16037 25143
rect 15988 25112 16037 25140
rect 15988 25100 15994 25112
rect 16025 25109 16037 25112
rect 16071 25109 16083 25143
rect 19794 25140 19800 25152
rect 19755 25112 19800 25140
rect 16025 25103 16083 25109
rect 19794 25100 19800 25112
rect 19852 25100 19858 25152
rect 22278 25100 22284 25152
rect 22336 25140 22342 25152
rect 23308 25149 23336 25248
rect 23661 25245 23673 25279
rect 23707 25276 23719 25279
rect 24486 25276 24492 25288
rect 23707 25248 24492 25276
rect 23707 25245 23719 25248
rect 23661 25239 23719 25245
rect 24486 25236 24492 25248
rect 24544 25236 24550 25288
rect 24946 25276 24952 25288
rect 24907 25248 24952 25276
rect 24946 25236 24952 25248
rect 25004 25236 25010 25288
rect 25777 25279 25835 25285
rect 25777 25245 25789 25279
rect 25823 25245 25835 25279
rect 25777 25239 25835 25245
rect 24670 25208 24676 25220
rect 24504 25180 24676 25208
rect 24504 25152 24532 25180
rect 24670 25168 24676 25180
rect 24728 25208 24734 25220
rect 25792 25208 25820 25239
rect 29362 25236 29368 25288
rect 29420 25276 29426 25288
rect 29730 25276 29736 25288
rect 29420 25248 29736 25276
rect 29420 25236 29426 25248
rect 29730 25236 29736 25248
rect 29788 25236 29794 25288
rect 30374 25276 30380 25288
rect 30335 25248 30380 25276
rect 30374 25236 30380 25248
rect 30432 25236 30438 25288
rect 30469 25279 30527 25285
rect 30469 25245 30481 25279
rect 30515 25245 30527 25279
rect 31386 25276 31392 25288
rect 31347 25248 31392 25276
rect 30469 25239 30527 25245
rect 26878 25208 26884 25220
rect 24728 25180 25820 25208
rect 26839 25180 26884 25208
rect 24728 25168 24734 25180
rect 26878 25168 26884 25180
rect 26936 25168 26942 25220
rect 29270 25208 29276 25220
rect 28106 25180 29276 25208
rect 29270 25168 29276 25180
rect 29328 25168 29334 25220
rect 30484 25208 30512 25239
rect 31386 25236 31392 25248
rect 31444 25236 31450 25288
rect 32217 25279 32275 25285
rect 32217 25245 32229 25279
rect 32263 25276 32275 25279
rect 33042 25276 33048 25288
rect 32263 25248 33048 25276
rect 32263 25245 32275 25248
rect 32217 25239 32275 25245
rect 33042 25236 33048 25248
rect 33100 25236 33106 25288
rect 34057 25279 34115 25285
rect 34057 25276 34069 25279
rect 33244 25248 34069 25276
rect 33244 25220 33272 25248
rect 34057 25245 34069 25248
rect 34103 25245 34115 25279
rect 34238 25276 34244 25288
rect 34199 25248 34244 25276
rect 34057 25239 34115 25245
rect 34238 25236 34244 25248
rect 34296 25236 34302 25288
rect 35084 25285 35112 25316
rect 35069 25279 35127 25285
rect 35069 25245 35081 25279
rect 35115 25245 35127 25279
rect 35069 25239 35127 25245
rect 35161 25279 35219 25285
rect 35161 25245 35173 25279
rect 35207 25245 35219 25279
rect 35161 25239 35219 25245
rect 30392 25180 30512 25208
rect 30392 25152 30420 25180
rect 32306 25168 32312 25220
rect 32364 25208 32370 25220
rect 32401 25211 32459 25217
rect 32401 25208 32413 25211
rect 32364 25180 32413 25208
rect 32364 25168 32370 25180
rect 32401 25177 32413 25180
rect 32447 25177 32459 25211
rect 33226 25208 33232 25220
rect 33187 25180 33232 25208
rect 32401 25171 32459 25177
rect 33226 25168 33232 25180
rect 33284 25168 33290 25220
rect 33413 25211 33471 25217
rect 33413 25177 33425 25211
rect 33459 25208 33471 25211
rect 33686 25208 33692 25220
rect 33459 25180 33692 25208
rect 33459 25177 33471 25180
rect 33413 25171 33471 25177
rect 33686 25168 33692 25180
rect 33744 25168 33750 25220
rect 34146 25208 34152 25220
rect 34059 25180 34152 25208
rect 34146 25168 34152 25180
rect 34204 25208 34210 25220
rect 35176 25208 35204 25239
rect 35526 25236 35532 25288
rect 35584 25276 35590 25288
rect 35713 25279 35771 25285
rect 35713 25276 35725 25279
rect 35584 25248 35725 25276
rect 35584 25236 35590 25248
rect 35713 25245 35725 25248
rect 35759 25245 35771 25279
rect 36354 25276 36360 25288
rect 36315 25248 36360 25276
rect 35713 25239 35771 25245
rect 36354 25236 36360 25248
rect 36412 25236 36418 25288
rect 34204 25180 35204 25208
rect 34204 25168 34210 25180
rect 22465 25143 22523 25149
rect 22465 25140 22477 25143
rect 22336 25112 22477 25140
rect 22336 25100 22342 25112
rect 22465 25109 22477 25112
rect 22511 25109 22523 25143
rect 22465 25103 22523 25109
rect 23293 25143 23351 25149
rect 23293 25109 23305 25143
rect 23339 25109 23351 25143
rect 23293 25103 23351 25109
rect 24486 25100 24492 25152
rect 24544 25100 24550 25152
rect 24854 25140 24860 25152
rect 24815 25112 24860 25140
rect 24854 25100 24860 25112
rect 24912 25100 24918 25152
rect 25317 25143 25375 25149
rect 25317 25109 25329 25143
rect 25363 25140 25375 25143
rect 25682 25140 25688 25152
rect 25363 25112 25688 25140
rect 25363 25109 25375 25112
rect 25317 25103 25375 25109
rect 25682 25100 25688 25112
rect 25740 25100 25746 25152
rect 25866 25140 25872 25152
rect 25827 25112 25872 25140
rect 25866 25100 25872 25112
rect 25924 25100 25930 25152
rect 30374 25100 30380 25152
rect 30432 25100 30438 25152
rect 33704 25140 33732 25168
rect 34238 25140 34244 25152
rect 33704 25112 34244 25140
rect 34238 25100 34244 25112
rect 34296 25100 34302 25152
rect 34790 25100 34796 25152
rect 34848 25140 34854 25152
rect 34885 25143 34943 25149
rect 34885 25140 34897 25143
rect 34848 25112 34897 25140
rect 34848 25100 34854 25112
rect 34885 25109 34897 25112
rect 34931 25109 34943 25143
rect 34885 25103 34943 25109
rect 1104 25050 37628 25072
rect 1104 24998 4874 25050
rect 4926 24998 4938 25050
rect 4990 24998 5002 25050
rect 5054 24998 5066 25050
rect 5118 24998 5130 25050
rect 5182 24998 35594 25050
rect 35646 24998 35658 25050
rect 35710 24998 35722 25050
rect 35774 24998 35786 25050
rect 35838 24998 35850 25050
rect 35902 24998 37628 25050
rect 1104 24976 37628 24998
rect 10686 24936 10692 24948
rect 10599 24908 10692 24936
rect 10686 24896 10692 24908
rect 10744 24936 10750 24948
rect 12066 24936 12072 24948
rect 10744 24908 12072 24936
rect 10744 24896 10750 24908
rect 12066 24896 12072 24908
rect 12124 24896 12130 24948
rect 21082 24936 21088 24948
rect 21043 24908 21088 24936
rect 21082 24896 21088 24908
rect 21140 24896 21146 24948
rect 23750 24936 23756 24948
rect 23711 24908 23756 24936
rect 23750 24896 23756 24908
rect 23808 24896 23814 24948
rect 24854 24896 24860 24948
rect 24912 24936 24918 24948
rect 25498 24936 25504 24948
rect 24912 24908 25504 24936
rect 24912 24896 24918 24908
rect 25498 24896 25504 24908
rect 25556 24936 25562 24948
rect 25961 24939 26019 24945
rect 25961 24936 25973 24939
rect 25556 24908 25973 24936
rect 25556 24896 25562 24908
rect 25961 24905 25973 24908
rect 26007 24905 26019 24939
rect 25961 24899 26019 24905
rect 26878 24896 26884 24948
rect 26936 24936 26942 24948
rect 27157 24939 27215 24945
rect 27157 24936 27169 24939
rect 26936 24908 27169 24936
rect 26936 24896 26942 24908
rect 27157 24905 27169 24908
rect 27203 24905 27215 24939
rect 27157 24899 27215 24905
rect 28902 24896 28908 24948
rect 28960 24936 28966 24948
rect 28997 24939 29055 24945
rect 28997 24936 29009 24939
rect 28960 24908 29009 24936
rect 28960 24896 28966 24908
rect 28997 24905 29009 24908
rect 29043 24905 29055 24939
rect 28997 24899 29055 24905
rect 30101 24939 30159 24945
rect 30101 24905 30113 24939
rect 30147 24936 30159 24939
rect 30282 24936 30288 24948
rect 30147 24908 30288 24936
rect 30147 24905 30159 24908
rect 30101 24899 30159 24905
rect 30282 24896 30288 24908
rect 30340 24896 30346 24948
rect 30558 24896 30564 24948
rect 30616 24936 30622 24948
rect 34790 24936 34796 24948
rect 30616 24908 31754 24936
rect 34751 24908 34796 24936
rect 30616 24896 30622 24908
rect 7742 24868 7748 24880
rect 7703 24840 7748 24868
rect 7742 24828 7748 24840
rect 7800 24828 7806 24880
rect 8478 24828 8484 24880
rect 8536 24828 8542 24880
rect 9674 24828 9680 24880
rect 9732 24868 9738 24880
rect 10134 24868 10140 24880
rect 9732 24840 10140 24868
rect 9732 24828 9738 24840
rect 10134 24828 10140 24840
rect 10192 24868 10198 24880
rect 10781 24871 10839 24877
rect 10781 24868 10793 24871
rect 10192 24840 10793 24868
rect 10192 24828 10198 24840
rect 10781 24837 10793 24840
rect 10827 24837 10839 24871
rect 10781 24831 10839 24837
rect 13265 24871 13323 24877
rect 13265 24837 13277 24871
rect 13311 24868 13323 24871
rect 14734 24868 14740 24880
rect 13311 24840 14740 24868
rect 13311 24837 13323 24840
rect 13265 24831 13323 24837
rect 14734 24828 14740 24840
rect 14792 24828 14798 24880
rect 19058 24868 19064 24880
rect 15212 24840 15608 24868
rect 19019 24840 19064 24868
rect 9769 24803 9827 24809
rect 9769 24800 9781 24803
rect 9508 24772 9781 24800
rect 7469 24735 7527 24741
rect 7469 24701 7481 24735
rect 7515 24701 7527 24735
rect 7469 24695 7527 24701
rect 7484 24596 7512 24695
rect 9508 24664 9536 24772
rect 9769 24769 9781 24772
rect 9815 24769 9827 24803
rect 9769 24763 9827 24769
rect 9861 24803 9919 24809
rect 9861 24769 9873 24803
rect 9907 24800 9919 24803
rect 9950 24800 9956 24812
rect 9907 24772 9956 24800
rect 9907 24769 9919 24772
rect 9861 24763 9919 24769
rect 9950 24760 9956 24772
rect 10008 24760 10014 24812
rect 11330 24760 11336 24812
rect 11388 24800 11394 24812
rect 14921 24803 14979 24809
rect 11388 24772 12388 24800
rect 11388 24760 11394 24772
rect 9582 24692 9588 24744
rect 9640 24732 9646 24744
rect 10505 24735 10563 24741
rect 10505 24732 10517 24735
rect 9640 24704 10517 24732
rect 9640 24692 9646 24704
rect 10505 24701 10517 24704
rect 10551 24701 10563 24735
rect 12158 24732 12164 24744
rect 12119 24704 12164 24732
rect 10505 24695 10563 24701
rect 12158 24692 12164 24704
rect 12216 24692 12222 24744
rect 12360 24741 12388 24772
rect 14921 24769 14933 24803
rect 14967 24800 14979 24803
rect 15212 24800 15240 24840
rect 14967 24772 15240 24800
rect 14967 24769 14979 24772
rect 14921 24763 14979 24769
rect 15286 24760 15292 24812
rect 15344 24800 15350 24812
rect 15580 24809 15608 24840
rect 19058 24828 19064 24840
rect 19116 24828 19122 24880
rect 20990 24868 20996 24880
rect 20951 24840 20996 24868
rect 20990 24828 20996 24840
rect 21048 24828 21054 24880
rect 22278 24868 22284 24880
rect 22239 24840 22284 24868
rect 22278 24828 22284 24840
rect 22336 24828 22342 24880
rect 25866 24868 25872 24880
rect 25714 24840 25872 24868
rect 25866 24828 25872 24840
rect 25924 24828 25930 24880
rect 29086 24868 29092 24880
rect 29047 24840 29092 24868
rect 29086 24828 29092 24840
rect 29144 24828 29150 24880
rect 30742 24868 30748 24880
rect 29196 24840 30748 24868
rect 15473 24803 15531 24809
rect 15473 24800 15485 24803
rect 15344 24772 15485 24800
rect 15344 24760 15350 24772
rect 15473 24769 15485 24772
rect 15519 24769 15531 24803
rect 15473 24763 15531 24769
rect 15565 24803 15623 24809
rect 15565 24769 15577 24803
rect 15611 24769 15623 24803
rect 15565 24763 15623 24769
rect 16117 24803 16175 24809
rect 16117 24769 16129 24803
rect 16163 24800 16175 24803
rect 17313 24803 17371 24809
rect 16163 24772 17264 24800
rect 16163 24769 16175 24772
rect 16117 24763 16175 24769
rect 12345 24735 12403 24741
rect 12345 24701 12357 24735
rect 12391 24732 12403 24735
rect 12986 24732 12992 24744
rect 12391 24704 12992 24732
rect 12391 24701 12403 24704
rect 12345 24695 12403 24701
rect 12986 24692 12992 24704
rect 13044 24692 13050 24744
rect 13170 24732 13176 24744
rect 13131 24704 13176 24732
rect 13170 24692 13176 24704
rect 13228 24692 13234 24744
rect 14829 24735 14887 24741
rect 14829 24701 14841 24735
rect 14875 24732 14887 24735
rect 15194 24732 15200 24744
rect 14875 24704 15200 24732
rect 14875 24701 14887 24704
rect 14829 24695 14887 24701
rect 15194 24692 15200 24704
rect 15252 24692 15258 24744
rect 15580 24732 15608 24763
rect 16758 24732 16764 24744
rect 15580 24704 16764 24732
rect 16758 24692 16764 24704
rect 16816 24692 16822 24744
rect 17037 24735 17095 24741
rect 17037 24701 17049 24735
rect 17083 24701 17095 24735
rect 17037 24695 17095 24701
rect 9858 24664 9864 24676
rect 9508 24636 9864 24664
rect 9858 24624 9864 24636
rect 9916 24664 9922 24676
rect 10870 24664 10876 24676
rect 9916 24636 10876 24664
rect 9916 24624 9922 24636
rect 10870 24624 10876 24636
rect 10928 24624 10934 24676
rect 10962 24624 10968 24676
rect 11020 24664 11026 24676
rect 11701 24667 11759 24673
rect 11701 24664 11713 24667
rect 11020 24636 11713 24664
rect 11020 24624 11026 24636
rect 11701 24633 11713 24636
rect 11747 24633 11759 24667
rect 11701 24627 11759 24633
rect 14458 24624 14464 24676
rect 14516 24664 14522 24676
rect 17052 24664 17080 24695
rect 14516 24636 17080 24664
rect 14516 24624 14522 24636
rect 9122 24596 9128 24608
rect 7484 24568 9128 24596
rect 9122 24556 9128 24568
rect 9180 24556 9186 24608
rect 9214 24556 9220 24608
rect 9272 24596 9278 24608
rect 9272 24568 9317 24596
rect 9272 24556 9278 24568
rect 10778 24556 10784 24608
rect 10836 24596 10842 24608
rect 11149 24599 11207 24605
rect 11149 24596 11161 24599
rect 10836 24568 11161 24596
rect 10836 24556 10842 24568
rect 11149 24565 11161 24568
rect 11195 24565 11207 24599
rect 11149 24559 11207 24565
rect 13538 24556 13544 24608
rect 13596 24596 13602 24608
rect 13633 24599 13691 24605
rect 13633 24596 13645 24599
rect 13596 24568 13645 24596
rect 13596 24556 13602 24568
rect 13633 24565 13645 24568
rect 13679 24565 13691 24599
rect 13633 24559 13691 24565
rect 16301 24599 16359 24605
rect 16301 24565 16313 24599
rect 16347 24596 16359 24599
rect 17126 24596 17132 24608
rect 16347 24568 17132 24596
rect 16347 24565 16359 24568
rect 16301 24559 16359 24565
rect 17126 24556 17132 24568
rect 17184 24556 17190 24608
rect 17236 24596 17264 24772
rect 17313 24769 17325 24803
rect 17359 24769 17371 24803
rect 17313 24763 17371 24769
rect 17328 24732 17356 24763
rect 17862 24760 17868 24812
rect 17920 24800 17926 24812
rect 17957 24803 18015 24809
rect 17957 24800 17969 24803
rect 17920 24772 17969 24800
rect 17920 24760 17926 24772
rect 17957 24769 17969 24772
rect 18003 24769 18015 24803
rect 17957 24763 18015 24769
rect 19153 24803 19211 24809
rect 19153 24769 19165 24803
rect 19199 24800 19211 24803
rect 19794 24800 19800 24812
rect 19199 24772 19800 24800
rect 19199 24769 19211 24772
rect 19153 24763 19211 24769
rect 19794 24760 19800 24772
rect 19852 24760 19858 24812
rect 20165 24803 20223 24809
rect 20165 24769 20177 24803
rect 20211 24800 20223 24803
rect 20346 24800 20352 24812
rect 20211 24772 20352 24800
rect 20211 24769 20223 24772
rect 20165 24763 20223 24769
rect 20346 24760 20352 24772
rect 20404 24760 20410 24812
rect 23658 24800 23664 24812
rect 23414 24772 23664 24800
rect 23658 24760 23664 24772
rect 23716 24760 23722 24812
rect 25774 24760 25780 24812
rect 25832 24800 25838 24812
rect 26605 24803 26663 24809
rect 26605 24800 26617 24803
rect 25832 24772 26617 24800
rect 25832 24760 25838 24772
rect 26605 24769 26617 24772
rect 26651 24769 26663 24803
rect 26605 24763 26663 24769
rect 27062 24760 27068 24812
rect 27120 24800 27126 24812
rect 27341 24803 27399 24809
rect 27341 24800 27353 24803
rect 27120 24772 27353 24800
rect 27120 24760 27126 24772
rect 27341 24769 27353 24772
rect 27387 24769 27399 24803
rect 27341 24763 27399 24769
rect 27430 24760 27436 24812
rect 27488 24800 27494 24812
rect 27801 24803 27859 24809
rect 27801 24800 27813 24803
rect 27488 24772 27813 24800
rect 27488 24760 27494 24772
rect 27801 24769 27813 24772
rect 27847 24769 27859 24803
rect 27801 24763 27859 24769
rect 27890 24760 27896 24812
rect 27948 24800 27954 24812
rect 28905 24803 28963 24809
rect 27948 24772 27993 24800
rect 27948 24760 27954 24772
rect 28905 24769 28917 24803
rect 28951 24800 28963 24803
rect 29196 24800 29224 24840
rect 30742 24828 30748 24840
rect 30800 24868 30806 24880
rect 31478 24868 31484 24880
rect 30800 24840 31484 24868
rect 30800 24828 30806 24840
rect 31478 24828 31484 24840
rect 31536 24828 31542 24880
rect 31726 24868 31754 24908
rect 34790 24896 34796 24908
rect 34848 24896 34854 24948
rect 31726 24840 33916 24868
rect 29730 24800 29736 24812
rect 28951 24772 29224 24800
rect 29691 24772 29736 24800
rect 28951 24769 28963 24772
rect 28905 24763 28963 24769
rect 29730 24760 29736 24772
rect 29788 24760 29794 24812
rect 30006 24760 30012 24812
rect 30064 24800 30070 24812
rect 30561 24803 30619 24809
rect 30561 24800 30573 24803
rect 30064 24772 30573 24800
rect 30064 24760 30070 24772
rect 30561 24769 30573 24772
rect 30607 24769 30619 24803
rect 30561 24763 30619 24769
rect 31202 24760 31208 24812
rect 31260 24800 31266 24812
rect 31297 24803 31355 24809
rect 31297 24800 31309 24803
rect 31260 24772 31309 24800
rect 31260 24760 31266 24772
rect 31297 24769 31309 24772
rect 31343 24769 31355 24803
rect 31297 24763 31355 24769
rect 31389 24803 31447 24809
rect 31389 24769 31401 24803
rect 31435 24769 31447 24803
rect 31389 24763 31447 24769
rect 18046 24732 18052 24744
rect 17328 24704 18052 24732
rect 18046 24692 18052 24704
rect 18104 24692 18110 24744
rect 18230 24692 18236 24744
rect 18288 24732 18294 24744
rect 18966 24732 18972 24744
rect 18288 24704 18972 24732
rect 18288 24692 18294 24704
rect 18966 24692 18972 24704
rect 19024 24732 19030 24744
rect 19245 24735 19303 24741
rect 19245 24732 19257 24735
rect 19024 24704 19257 24732
rect 19024 24692 19030 24704
rect 19245 24701 19257 24704
rect 19291 24701 19303 24735
rect 19245 24695 19303 24701
rect 20806 24692 20812 24744
rect 20864 24732 20870 24744
rect 21269 24735 21327 24741
rect 21269 24732 21281 24735
rect 20864 24704 21281 24732
rect 20864 24692 20870 24704
rect 21269 24701 21281 24704
rect 21315 24732 21327 24735
rect 21818 24732 21824 24744
rect 21315 24704 21824 24732
rect 21315 24701 21327 24704
rect 21269 24695 21327 24701
rect 21818 24692 21824 24704
rect 21876 24692 21882 24744
rect 22005 24735 22063 24741
rect 22005 24701 22017 24735
rect 22051 24701 22063 24735
rect 22005 24695 22063 24701
rect 24213 24735 24271 24741
rect 24213 24701 24225 24735
rect 24259 24701 24271 24735
rect 24213 24695 24271 24701
rect 24489 24735 24547 24741
rect 24489 24701 24501 24735
rect 24535 24732 24547 24735
rect 24535 24704 25544 24732
rect 24535 24701 24547 24704
rect 24489 24695 24547 24701
rect 17865 24667 17923 24673
rect 17865 24633 17877 24667
rect 17911 24664 17923 24667
rect 17954 24664 17960 24676
rect 17911 24636 17960 24664
rect 17911 24633 17923 24636
rect 17865 24627 17923 24633
rect 17954 24624 17960 24636
rect 18012 24624 18018 24676
rect 20625 24667 20683 24673
rect 20625 24664 20637 24667
rect 18064 24636 20637 24664
rect 18064 24596 18092 24636
rect 20625 24633 20637 24636
rect 20671 24633 20683 24667
rect 20625 24627 20683 24633
rect 17236 24568 18092 24596
rect 18322 24556 18328 24608
rect 18380 24596 18386 24608
rect 18693 24599 18751 24605
rect 18693 24596 18705 24599
rect 18380 24568 18705 24596
rect 18380 24556 18386 24568
rect 18693 24565 18705 24568
rect 18739 24565 18751 24599
rect 19978 24596 19984 24608
rect 19939 24568 19984 24596
rect 18693 24559 18751 24565
rect 19978 24556 19984 24568
rect 20036 24556 20042 24608
rect 22020 24596 22048 24695
rect 22738 24596 22744 24608
rect 22020 24568 22744 24596
rect 22738 24556 22744 24568
rect 22796 24596 22802 24608
rect 24228 24596 24256 24695
rect 25516 24664 25544 24704
rect 29454 24692 29460 24744
rect 29512 24732 29518 24744
rect 29825 24735 29883 24741
rect 29825 24732 29837 24735
rect 29512 24704 29837 24732
rect 29512 24692 29518 24704
rect 29825 24701 29837 24704
rect 29871 24701 29883 24735
rect 29825 24695 29883 24701
rect 29914 24692 29920 24744
rect 29972 24732 29978 24744
rect 30650 24732 30656 24744
rect 29972 24704 30656 24732
rect 29972 24692 29978 24704
rect 30650 24692 30656 24704
rect 30708 24692 30714 24744
rect 31404 24676 31432 24763
rect 32490 24760 32496 24812
rect 32548 24800 32554 24812
rect 32769 24803 32827 24809
rect 32769 24800 32781 24803
rect 32548 24772 32781 24800
rect 32548 24760 32554 24772
rect 32769 24769 32781 24772
rect 32815 24769 32827 24803
rect 32769 24763 32827 24769
rect 32953 24803 33011 24809
rect 32953 24769 32965 24803
rect 32999 24769 33011 24803
rect 32953 24763 33011 24769
rect 32214 24692 32220 24744
rect 32272 24732 32278 24744
rect 32968 24732 32996 24763
rect 33226 24760 33232 24812
rect 33284 24800 33290 24812
rect 33781 24803 33839 24809
rect 33781 24800 33793 24803
rect 33284 24772 33793 24800
rect 33284 24760 33290 24772
rect 33781 24769 33793 24772
rect 33827 24769 33839 24803
rect 33888 24800 33916 24840
rect 36354 24800 36360 24812
rect 33888 24772 34560 24800
rect 33781 24763 33839 24769
rect 32272 24704 32996 24732
rect 32272 24692 32278 24704
rect 33502 24692 33508 24744
rect 33560 24732 33566 24744
rect 34532 24741 34560 24772
rect 35866 24772 36360 24800
rect 33597 24735 33655 24741
rect 33597 24732 33609 24735
rect 33560 24704 33609 24732
rect 33560 24692 33566 24704
rect 33597 24701 33609 24704
rect 33643 24701 33655 24735
rect 33597 24695 33655 24701
rect 34517 24735 34575 24741
rect 34517 24701 34529 24735
rect 34563 24701 34575 24735
rect 34698 24732 34704 24744
rect 34659 24704 34704 24732
rect 34517 24695 34575 24701
rect 26421 24667 26479 24673
rect 26421 24664 26433 24667
rect 25516 24636 26433 24664
rect 26421 24633 26433 24636
rect 26467 24633 26479 24667
rect 26421 24627 26479 24633
rect 28721 24667 28779 24673
rect 28721 24633 28733 24667
rect 28767 24633 28779 24667
rect 28721 24627 28779 24633
rect 29273 24667 29331 24673
rect 29273 24633 29285 24667
rect 29319 24664 29331 24667
rect 30466 24664 30472 24676
rect 29319 24636 30472 24664
rect 29319 24633 29331 24636
rect 29273 24627 29331 24633
rect 27154 24596 27160 24608
rect 22796 24568 27160 24596
rect 22796 24556 22802 24568
rect 27154 24556 27160 24568
rect 27212 24556 27218 24608
rect 28736 24596 28764 24627
rect 30466 24624 30472 24636
rect 30524 24624 30530 24676
rect 31386 24624 31392 24676
rect 31444 24664 31450 24676
rect 34532 24664 34560 24695
rect 34698 24692 34704 24704
rect 34756 24692 34762 24744
rect 34606 24664 34612 24676
rect 31444 24636 34100 24664
rect 34532 24636 34612 24664
rect 31444 24624 31450 24636
rect 28994 24596 29000 24608
rect 28736 24568 29000 24596
rect 28994 24556 29000 24568
rect 29052 24596 29058 24608
rect 29822 24596 29828 24608
rect 29052 24568 29828 24596
rect 29052 24556 29058 24568
rect 29822 24556 29828 24568
rect 29880 24556 29886 24608
rect 29917 24599 29975 24605
rect 29917 24565 29929 24599
rect 29963 24596 29975 24599
rect 30006 24596 30012 24608
rect 29963 24568 30012 24596
rect 29963 24565 29975 24568
rect 29917 24559 29975 24565
rect 30006 24556 30012 24568
rect 30064 24556 30070 24608
rect 30374 24556 30380 24608
rect 30432 24596 30438 24608
rect 30653 24599 30711 24605
rect 30653 24596 30665 24599
rect 30432 24568 30665 24596
rect 30432 24556 30438 24568
rect 30653 24565 30665 24568
rect 30699 24565 30711 24599
rect 30653 24559 30711 24565
rect 33137 24599 33195 24605
rect 33137 24565 33149 24599
rect 33183 24596 33195 24599
rect 33778 24596 33784 24608
rect 33183 24568 33784 24596
rect 33183 24565 33195 24568
rect 33137 24559 33195 24565
rect 33778 24556 33784 24568
rect 33836 24556 33842 24608
rect 33962 24596 33968 24608
rect 33923 24568 33968 24596
rect 33962 24556 33968 24568
rect 34020 24556 34026 24608
rect 34072 24596 34100 24636
rect 34606 24624 34612 24636
rect 34664 24624 34670 24676
rect 35866 24664 35894 24772
rect 36354 24760 36360 24772
rect 36412 24760 36418 24812
rect 36446 24760 36452 24812
rect 36504 24800 36510 24812
rect 36504 24772 36549 24800
rect 36504 24760 36510 24772
rect 34716 24636 35894 24664
rect 34716 24596 34744 24636
rect 34072 24568 34744 24596
rect 35161 24599 35219 24605
rect 35161 24565 35173 24599
rect 35207 24596 35219 24599
rect 35342 24596 35348 24608
rect 35207 24568 35348 24596
rect 35207 24565 35219 24568
rect 35161 24559 35219 24565
rect 35342 24556 35348 24568
rect 35400 24556 35406 24608
rect 1104 24506 37628 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 37628 24506
rect 1104 24432 37628 24454
rect 7837 24395 7895 24401
rect 7837 24361 7849 24395
rect 7883 24392 7895 24395
rect 7926 24392 7932 24404
rect 7883 24364 7932 24392
rect 7883 24361 7895 24364
rect 7837 24355 7895 24361
rect 7926 24352 7932 24364
rect 7984 24352 7990 24404
rect 15654 24392 15660 24404
rect 15615 24364 15660 24392
rect 15654 24352 15660 24364
rect 15712 24352 15718 24404
rect 16942 24352 16948 24404
rect 17000 24392 17006 24404
rect 20346 24392 20352 24404
rect 17000 24364 17448 24392
rect 20307 24364 20352 24392
rect 17000 24352 17006 24364
rect 8110 24284 8116 24336
rect 8168 24324 8174 24336
rect 11330 24324 11336 24336
rect 8168 24296 11336 24324
rect 8168 24284 8174 24296
rect 8202 24216 8208 24268
rect 8260 24256 8266 24268
rect 8496 24265 8524 24296
rect 11330 24284 11336 24296
rect 11388 24284 11394 24336
rect 8297 24259 8355 24265
rect 8297 24256 8309 24259
rect 8260 24228 8309 24256
rect 8260 24216 8266 24228
rect 8297 24225 8309 24228
rect 8343 24225 8355 24259
rect 8297 24219 8355 24225
rect 8481 24259 8539 24265
rect 8481 24225 8493 24259
rect 8527 24225 8539 24259
rect 8481 24219 8539 24225
rect 9122 24216 9128 24268
rect 9180 24256 9186 24268
rect 9766 24256 9772 24268
rect 9180 24228 9772 24256
rect 9180 24216 9186 24228
rect 9766 24216 9772 24228
rect 9824 24256 9830 24268
rect 10045 24259 10103 24265
rect 10045 24256 10057 24259
rect 9824 24228 10057 24256
rect 9824 24216 9830 24228
rect 10045 24225 10057 24228
rect 10091 24225 10103 24259
rect 10045 24219 10103 24225
rect 11146 24216 11152 24268
rect 11204 24256 11210 24268
rect 11698 24256 11704 24268
rect 11204 24228 11704 24256
rect 11204 24216 11210 24228
rect 11698 24216 11704 24228
rect 11756 24256 11762 24268
rect 12342 24256 12348 24268
rect 11756 24228 12348 24256
rect 11756 24216 11762 24228
rect 12342 24216 12348 24228
rect 12400 24256 12406 24268
rect 12713 24259 12771 24265
rect 12713 24256 12725 24259
rect 12400 24228 12725 24256
rect 12400 24216 12406 24228
rect 12713 24225 12725 24228
rect 12759 24225 12771 24259
rect 17126 24256 17132 24268
rect 17087 24228 17132 24256
rect 12713 24219 12771 24225
rect 17126 24216 17132 24228
rect 17184 24216 17190 24268
rect 17420 24265 17448 24364
rect 20346 24352 20352 24364
rect 20404 24352 20410 24404
rect 23658 24392 23664 24404
rect 23619 24364 23664 24392
rect 23658 24352 23664 24364
rect 23716 24352 23722 24404
rect 27062 24392 27068 24404
rect 27023 24364 27068 24392
rect 27062 24352 27068 24364
rect 27120 24352 27126 24404
rect 30466 24392 30472 24404
rect 29012 24364 30472 24392
rect 17862 24284 17868 24336
rect 17920 24324 17926 24336
rect 29012 24324 29040 24364
rect 30466 24352 30472 24364
rect 30524 24352 30530 24404
rect 17920 24296 29040 24324
rect 17920 24284 17926 24296
rect 17405 24259 17463 24265
rect 17405 24225 17417 24259
rect 17451 24256 17463 24259
rect 17451 24228 18460 24256
rect 17451 24225 17463 24228
rect 17405 24219 17463 24225
rect 1765 24191 1823 24197
rect 1765 24157 1777 24191
rect 1811 24188 1823 24191
rect 2222 24188 2228 24200
rect 1811 24160 2228 24188
rect 1811 24157 1823 24160
rect 1765 24151 1823 24157
rect 2222 24148 2228 24160
rect 2280 24148 2286 24200
rect 7377 24191 7435 24197
rect 7377 24157 7389 24191
rect 7423 24188 7435 24191
rect 9858 24188 9864 24200
rect 7423 24160 9864 24188
rect 7423 24157 7435 24160
rect 7377 24151 7435 24157
rect 9858 24148 9864 24160
rect 9916 24148 9922 24200
rect 11330 24188 11336 24200
rect 11291 24160 11336 24188
rect 11330 24148 11336 24160
rect 11388 24148 11394 24200
rect 13538 24188 13544 24200
rect 13499 24160 13544 24188
rect 13538 24148 13544 24160
rect 13596 24148 13602 24200
rect 14458 24188 14464 24200
rect 14419 24160 14464 24188
rect 14458 24148 14464 24160
rect 14516 24148 14522 24200
rect 15013 24191 15071 24197
rect 15013 24157 15025 24191
rect 15059 24157 15071 24191
rect 18322 24188 18328 24200
rect 18283 24160 18328 24188
rect 15013 24151 15071 24157
rect 8205 24123 8263 24129
rect 8205 24089 8217 24123
rect 8251 24120 8263 24123
rect 9214 24120 9220 24132
rect 8251 24092 9220 24120
rect 8251 24089 8263 24092
rect 8205 24083 8263 24089
rect 9214 24080 9220 24092
rect 9272 24080 9278 24132
rect 10873 24123 10931 24129
rect 10873 24089 10885 24123
rect 10919 24120 10931 24123
rect 11974 24120 11980 24132
rect 10919 24092 11980 24120
rect 10919 24089 10931 24092
rect 10873 24083 10931 24089
rect 11974 24080 11980 24092
rect 12032 24080 12038 24132
rect 15028 24120 15056 24151
rect 18322 24148 18328 24160
rect 18380 24148 18386 24200
rect 18432 24188 18460 24228
rect 19610 24216 19616 24268
rect 19668 24256 19674 24268
rect 19705 24259 19763 24265
rect 19705 24256 19717 24259
rect 19668 24228 19717 24256
rect 19668 24216 19674 24228
rect 19705 24225 19717 24228
rect 19751 24225 19763 24259
rect 19705 24219 19763 24225
rect 19794 24216 19800 24268
rect 19852 24256 19858 24268
rect 19889 24259 19947 24265
rect 19889 24256 19901 24259
rect 19852 24228 19901 24256
rect 19852 24216 19858 24228
rect 19889 24225 19901 24228
rect 19935 24225 19947 24259
rect 19889 24219 19947 24225
rect 19996 24228 22094 24256
rect 18598 24188 18604 24200
rect 18432 24160 18604 24188
rect 18598 24148 18604 24160
rect 18656 24188 18662 24200
rect 19996 24188 20024 24228
rect 18656 24160 20024 24188
rect 18656 24148 18662 24160
rect 20714 24148 20720 24200
rect 20772 24188 20778 24200
rect 21174 24188 21180 24200
rect 20772 24160 21180 24188
rect 20772 24148 20778 24160
rect 21174 24148 21180 24160
rect 21232 24188 21238 24200
rect 21269 24191 21327 24197
rect 21269 24188 21281 24191
rect 21232 24160 21281 24188
rect 21232 24148 21238 24160
rect 21269 24157 21281 24160
rect 21315 24157 21327 24191
rect 21269 24151 21327 24157
rect 15028 24092 15884 24120
rect 1578 24052 1584 24064
rect 1539 24024 1584 24052
rect 1578 24012 1584 24024
rect 1636 24012 1642 24064
rect 7282 24052 7288 24064
rect 7243 24024 7288 24052
rect 7282 24012 7288 24024
rect 7340 24012 7346 24064
rect 11517 24055 11575 24061
rect 11517 24021 11529 24055
rect 11563 24052 11575 24055
rect 11882 24052 11888 24064
rect 11563 24024 11888 24052
rect 11563 24021 11575 24024
rect 11517 24015 11575 24021
rect 11882 24012 11888 24024
rect 11940 24012 11946 24064
rect 13262 24012 13268 24064
rect 13320 24052 13326 24064
rect 13357 24055 13415 24061
rect 13357 24052 13369 24055
rect 13320 24024 13369 24052
rect 13320 24012 13326 24024
rect 13357 24021 13369 24024
rect 13403 24021 13415 24055
rect 14366 24052 14372 24064
rect 14327 24024 14372 24052
rect 13357 24015 13415 24021
rect 14366 24012 14372 24024
rect 14424 24012 14430 24064
rect 15197 24055 15255 24061
rect 15197 24021 15209 24055
rect 15243 24052 15255 24055
rect 15470 24052 15476 24064
rect 15243 24024 15476 24052
rect 15243 24021 15255 24024
rect 15197 24015 15255 24021
rect 15470 24012 15476 24024
rect 15528 24012 15534 24064
rect 15856 24052 15884 24092
rect 16666 24080 16672 24132
rect 16724 24080 16730 24132
rect 20898 24120 20904 24132
rect 17696 24092 20904 24120
rect 17696 24052 17724 24092
rect 20898 24080 20904 24092
rect 20956 24080 20962 24132
rect 22066 24120 22094 24228
rect 25590 24216 25596 24268
rect 25648 24256 25654 24268
rect 25685 24259 25743 24265
rect 25685 24256 25697 24259
rect 25648 24228 25697 24256
rect 25648 24216 25654 24228
rect 25685 24225 25697 24228
rect 25731 24225 25743 24259
rect 25685 24219 25743 24225
rect 25866 24216 25872 24268
rect 25924 24256 25930 24268
rect 26234 24256 26240 24268
rect 25924 24228 26240 24256
rect 25924 24216 25930 24228
rect 26234 24216 26240 24228
rect 26292 24256 26298 24268
rect 26421 24259 26479 24265
rect 26421 24256 26433 24259
rect 26292 24228 26433 24256
rect 26292 24216 26298 24228
rect 26421 24225 26433 24228
rect 26467 24225 26479 24259
rect 26421 24219 26479 24225
rect 23106 24188 23112 24200
rect 23067 24160 23112 24188
rect 23106 24148 23112 24160
rect 23164 24148 23170 24200
rect 23753 24191 23811 24197
rect 23753 24157 23765 24191
rect 23799 24188 23811 24191
rect 24486 24188 24492 24200
rect 23799 24160 24492 24188
rect 23799 24157 23811 24160
rect 23753 24151 23811 24157
rect 24486 24148 24492 24160
rect 24544 24148 24550 24200
rect 25498 24188 25504 24200
rect 25459 24160 25504 24188
rect 25498 24148 25504 24160
rect 25556 24188 25562 24200
rect 26605 24191 26663 24197
rect 26605 24188 26617 24191
rect 25556 24160 26617 24188
rect 25556 24148 25562 24160
rect 26605 24157 26617 24160
rect 26651 24157 26663 24191
rect 26605 24151 26663 24157
rect 26697 24191 26755 24197
rect 26697 24157 26709 24191
rect 26743 24188 26755 24191
rect 28350 24188 28356 24200
rect 26743 24160 28356 24188
rect 26743 24157 26755 24160
rect 26697 24151 26755 24157
rect 28350 24148 28356 24160
rect 28408 24148 28414 24200
rect 29012 24197 29040 24296
rect 32769 24327 32827 24333
rect 32769 24293 32781 24327
rect 32815 24324 32827 24327
rect 33502 24324 33508 24336
rect 32815 24296 33508 24324
rect 32815 24293 32827 24296
rect 32769 24287 32827 24293
rect 33502 24284 33508 24296
rect 33560 24284 33566 24336
rect 34698 24324 34704 24336
rect 33796 24296 34704 24324
rect 30466 24216 30472 24268
rect 30524 24256 30530 24268
rect 31481 24259 31539 24265
rect 31481 24256 31493 24259
rect 30524 24228 31493 24256
rect 30524 24216 30530 24228
rect 31481 24225 31493 24228
rect 31527 24225 31539 24259
rect 31481 24219 31539 24225
rect 31757 24259 31815 24265
rect 31757 24225 31769 24259
rect 31803 24256 31815 24259
rect 31938 24256 31944 24268
rect 31803 24228 31944 24256
rect 31803 24225 31815 24228
rect 31757 24219 31815 24225
rect 31938 24216 31944 24228
rect 31996 24216 32002 24268
rect 32030 24216 32036 24268
rect 32088 24256 32094 24268
rect 32306 24256 32312 24268
rect 32088 24228 32312 24256
rect 32088 24216 32094 24228
rect 32306 24216 32312 24228
rect 32364 24216 32370 24268
rect 32490 24216 32496 24268
rect 32548 24256 32554 24268
rect 33796 24265 33824 24296
rect 34698 24284 34704 24296
rect 34756 24284 34762 24336
rect 33781 24259 33839 24265
rect 33781 24256 33793 24259
rect 32548 24228 33793 24256
rect 32548 24216 32554 24228
rect 33781 24225 33793 24228
rect 33827 24225 33839 24259
rect 34146 24256 34152 24268
rect 34107 24228 34152 24256
rect 33781 24219 33839 24225
rect 34146 24216 34152 24228
rect 34204 24216 34210 24268
rect 34606 24216 34612 24268
rect 34664 24256 34670 24268
rect 35437 24259 35495 24265
rect 35437 24256 35449 24259
rect 34664 24228 35449 24256
rect 34664 24216 34670 24228
rect 35437 24225 35449 24228
rect 35483 24225 35495 24259
rect 35437 24219 35495 24225
rect 28997 24191 29055 24197
rect 28997 24157 29009 24191
rect 29043 24157 29055 24191
rect 28997 24151 29055 24157
rect 29089 24191 29147 24197
rect 29089 24157 29101 24191
rect 29135 24188 29147 24191
rect 29135 24160 30406 24188
rect 29135 24157 29147 24160
rect 29089 24151 29147 24157
rect 32214 24148 32220 24200
rect 32272 24188 32278 24200
rect 32401 24191 32459 24197
rect 32401 24188 32413 24191
rect 32272 24160 32413 24188
rect 32272 24148 32278 24160
rect 32401 24157 32413 24160
rect 32447 24157 32459 24191
rect 32401 24151 32459 24157
rect 29733 24123 29791 24129
rect 29733 24120 29745 24123
rect 22066 24092 29745 24120
rect 29733 24089 29745 24092
rect 29779 24089 29791 24123
rect 32416 24120 32444 24151
rect 33134 24148 33140 24200
rect 33192 24188 33198 24200
rect 33689 24191 33747 24197
rect 33689 24188 33701 24191
rect 33192 24160 33701 24188
rect 33192 24148 33198 24160
rect 33689 24157 33701 24160
rect 33735 24157 33747 24191
rect 36906 24188 36912 24200
rect 36867 24160 36912 24188
rect 33689 24151 33747 24157
rect 36906 24148 36912 24160
rect 36964 24148 36970 24200
rect 35345 24123 35403 24129
rect 35345 24120 35357 24123
rect 32416 24092 35357 24120
rect 29733 24083 29791 24089
rect 35345 24089 35357 24092
rect 35391 24120 35403 24123
rect 36814 24120 36820 24132
rect 35391 24092 36820 24120
rect 35391 24089 35403 24092
rect 35345 24083 35403 24089
rect 36814 24080 36820 24092
rect 36872 24080 36878 24132
rect 15856 24024 17724 24052
rect 17770 24012 17776 24064
rect 17828 24052 17834 24064
rect 18141 24055 18199 24061
rect 18141 24052 18153 24055
rect 17828 24024 18153 24052
rect 17828 24012 17834 24024
rect 18141 24021 18153 24024
rect 18187 24021 18199 24055
rect 18141 24015 18199 24021
rect 19886 24012 19892 24064
rect 19944 24052 19950 24064
rect 19981 24055 20039 24061
rect 19981 24052 19993 24055
rect 19944 24024 19993 24052
rect 19944 24012 19950 24024
rect 19981 24021 19993 24024
rect 20027 24021 20039 24055
rect 19981 24015 20039 24021
rect 21082 24012 21088 24064
rect 21140 24052 21146 24064
rect 21177 24055 21235 24061
rect 21177 24052 21189 24055
rect 21140 24024 21189 24052
rect 21140 24012 21146 24024
rect 21177 24021 21189 24024
rect 21223 24021 21235 24055
rect 21177 24015 21235 24021
rect 22554 24012 22560 24064
rect 22612 24052 22618 24064
rect 22925 24055 22983 24061
rect 22925 24052 22937 24055
rect 22612 24024 22937 24052
rect 22612 24012 22618 24024
rect 22925 24021 22937 24024
rect 22971 24021 22983 24055
rect 22925 24015 22983 24021
rect 24394 24012 24400 24064
rect 24452 24052 24458 24064
rect 25133 24055 25191 24061
rect 25133 24052 25145 24055
rect 24452 24024 25145 24052
rect 24452 24012 24458 24024
rect 25133 24021 25145 24024
rect 25179 24021 25191 24055
rect 25133 24015 25191 24021
rect 25593 24055 25651 24061
rect 25593 24021 25605 24055
rect 25639 24052 25651 24055
rect 26142 24052 26148 24064
rect 25639 24024 26148 24052
rect 25639 24021 25651 24024
rect 25593 24015 25651 24021
rect 26142 24012 26148 24024
rect 26200 24012 26206 24064
rect 33505 24055 33563 24061
rect 33505 24021 33517 24055
rect 33551 24052 33563 24055
rect 33594 24052 33600 24064
rect 33551 24024 33600 24052
rect 33551 24021 33563 24024
rect 33505 24015 33563 24021
rect 33594 24012 33600 24024
rect 33652 24012 33658 24064
rect 34422 24012 34428 24064
rect 34480 24052 34486 24064
rect 34885 24055 34943 24061
rect 34885 24052 34897 24055
rect 34480 24024 34897 24052
rect 34480 24012 34486 24024
rect 34885 24021 34897 24024
rect 34931 24021 34943 24055
rect 34885 24015 34943 24021
rect 34974 24012 34980 24064
rect 35032 24052 35038 24064
rect 35253 24055 35311 24061
rect 35253 24052 35265 24055
rect 35032 24024 35265 24052
rect 35032 24012 35038 24024
rect 35253 24021 35265 24024
rect 35299 24021 35311 24055
rect 37090 24052 37096 24064
rect 37051 24024 37096 24052
rect 35253 24015 35311 24021
rect 37090 24012 37096 24024
rect 37148 24012 37154 24064
rect 1104 23962 37628 23984
rect 1104 23910 4874 23962
rect 4926 23910 4938 23962
rect 4990 23910 5002 23962
rect 5054 23910 5066 23962
rect 5118 23910 5130 23962
rect 5182 23910 35594 23962
rect 35646 23910 35658 23962
rect 35710 23910 35722 23962
rect 35774 23910 35786 23962
rect 35838 23910 35850 23962
rect 35902 23910 37628 23962
rect 1104 23888 37628 23910
rect 9306 23808 9312 23860
rect 9364 23848 9370 23860
rect 9585 23851 9643 23857
rect 9585 23848 9597 23851
rect 9364 23820 9597 23848
rect 9364 23808 9370 23820
rect 9585 23817 9597 23820
rect 9631 23817 9643 23851
rect 10778 23848 10784 23860
rect 10739 23820 10784 23848
rect 9585 23811 9643 23817
rect 10778 23808 10784 23820
rect 10836 23808 10842 23860
rect 10873 23851 10931 23857
rect 10873 23817 10885 23851
rect 10919 23848 10931 23851
rect 12158 23848 12164 23860
rect 10919 23820 12164 23848
rect 10919 23817 10931 23820
rect 10873 23811 10931 23817
rect 12158 23808 12164 23820
rect 12216 23808 12222 23860
rect 14734 23848 14740 23860
rect 12406 23820 14740 23848
rect 7282 23740 7288 23792
rect 7340 23780 7346 23792
rect 7340 23752 7774 23780
rect 7340 23740 7346 23752
rect 10226 23740 10232 23792
rect 10284 23780 10290 23792
rect 12069 23783 12127 23789
rect 12069 23780 12081 23783
rect 10284 23752 12081 23780
rect 10284 23740 10290 23752
rect 12069 23749 12081 23752
rect 12115 23780 12127 23783
rect 12406 23780 12434 23820
rect 14734 23808 14740 23820
rect 14792 23848 14798 23860
rect 16574 23848 16580 23860
rect 14792 23820 16580 23848
rect 14792 23808 14798 23820
rect 16574 23808 16580 23820
rect 16632 23808 16638 23860
rect 16666 23808 16672 23860
rect 16724 23848 16730 23860
rect 16945 23851 17003 23857
rect 16945 23848 16957 23851
rect 16724 23820 16957 23848
rect 16724 23808 16730 23820
rect 16945 23817 16957 23820
rect 16991 23817 17003 23851
rect 17862 23848 17868 23860
rect 16945 23811 17003 23817
rect 17328 23820 17868 23848
rect 13262 23780 13268 23792
rect 12115 23752 12434 23780
rect 13223 23752 13268 23780
rect 12115 23749 12127 23752
rect 12069 23743 12127 23749
rect 13262 23740 13268 23752
rect 13320 23740 13326 23792
rect 8772 23684 12112 23712
rect 8772 23656 8800 23684
rect 6914 23604 6920 23656
rect 6972 23644 6978 23656
rect 7009 23647 7067 23653
rect 7009 23644 7021 23647
rect 6972 23616 7021 23644
rect 6972 23604 6978 23616
rect 7009 23613 7021 23616
rect 7055 23613 7067 23647
rect 7282 23644 7288 23656
rect 7243 23616 7288 23644
rect 7009 23607 7067 23613
rect 7282 23604 7288 23616
rect 7340 23604 7346 23656
rect 8754 23644 8760 23656
rect 8667 23616 8760 23644
rect 8754 23604 8760 23616
rect 8812 23604 8818 23656
rect 9674 23644 9680 23656
rect 9635 23616 9680 23644
rect 9674 23604 9680 23616
rect 9732 23604 9738 23656
rect 9766 23604 9772 23656
rect 9824 23644 9830 23656
rect 10965 23647 11023 23653
rect 10965 23644 10977 23647
rect 9824 23616 10977 23644
rect 9824 23604 9830 23616
rect 10965 23613 10977 23616
rect 11011 23644 11023 23647
rect 11790 23644 11796 23656
rect 11011 23616 11796 23644
rect 11011 23613 11023 23616
rect 10965 23607 11023 23613
rect 11790 23604 11796 23616
rect 11848 23604 11854 23656
rect 11977 23647 12035 23653
rect 11977 23613 11989 23647
rect 12023 23613 12035 23647
rect 12084 23644 12112 23684
rect 12342 23672 12348 23724
rect 12400 23712 12406 23724
rect 12989 23715 13047 23721
rect 12989 23712 13001 23715
rect 12400 23684 13001 23712
rect 12400 23672 12406 23684
rect 12989 23681 13001 23684
rect 13035 23681 13047 23715
rect 12989 23675 13047 23681
rect 14366 23672 14372 23724
rect 14424 23672 14430 23724
rect 15194 23672 15200 23724
rect 15252 23712 15258 23724
rect 15381 23715 15439 23721
rect 15381 23712 15393 23715
rect 15252 23684 15393 23712
rect 15252 23672 15258 23684
rect 15381 23681 15393 23684
rect 15427 23681 15439 23715
rect 15381 23675 15439 23681
rect 16758 23672 16764 23724
rect 16816 23712 16822 23724
rect 17037 23715 17095 23721
rect 17037 23712 17049 23715
rect 16816 23684 17049 23712
rect 16816 23672 16822 23684
rect 17037 23681 17049 23684
rect 17083 23712 17095 23715
rect 17328 23712 17356 23820
rect 17862 23808 17868 23820
rect 17920 23808 17926 23860
rect 19245 23851 19303 23857
rect 19245 23817 19257 23851
rect 19291 23848 19303 23851
rect 19794 23848 19800 23860
rect 19291 23820 19800 23848
rect 19291 23817 19303 23820
rect 19245 23811 19303 23817
rect 19794 23808 19800 23820
rect 19852 23808 19858 23860
rect 20806 23808 20812 23860
rect 20864 23848 20870 23860
rect 20864 23820 22094 23848
rect 20864 23808 20870 23820
rect 17770 23780 17776 23792
rect 17731 23752 17776 23780
rect 17770 23740 17776 23752
rect 17828 23740 17834 23792
rect 18506 23740 18512 23792
rect 18564 23740 18570 23792
rect 19978 23780 19984 23792
rect 19939 23752 19984 23780
rect 19978 23740 19984 23752
rect 20036 23740 20042 23792
rect 17083 23684 17356 23712
rect 17083 23681 17095 23684
rect 17037 23675 17095 23681
rect 21082 23672 21088 23724
rect 21140 23672 21146 23724
rect 22066 23712 22094 23820
rect 23106 23808 23112 23860
rect 23164 23848 23170 23860
rect 24029 23851 24087 23857
rect 24029 23848 24041 23851
rect 23164 23820 24041 23848
rect 23164 23808 23170 23820
rect 24029 23817 24041 23820
rect 24075 23817 24087 23851
rect 24394 23848 24400 23860
rect 24355 23820 24400 23848
rect 24029 23811 24087 23817
rect 24394 23808 24400 23820
rect 24452 23808 24458 23860
rect 26142 23848 26148 23860
rect 26055 23820 26148 23848
rect 26142 23808 26148 23820
rect 26200 23848 26206 23860
rect 28074 23848 28080 23860
rect 26200 23820 28080 23848
rect 26200 23808 26206 23820
rect 28074 23808 28080 23820
rect 28132 23848 28138 23860
rect 28905 23851 28963 23857
rect 28905 23848 28917 23851
rect 28132 23820 28917 23848
rect 28132 23808 28138 23820
rect 28905 23817 28917 23820
rect 28951 23817 28963 23851
rect 28905 23811 28963 23817
rect 32861 23851 32919 23857
rect 32861 23817 32873 23851
rect 32907 23848 32919 23851
rect 33226 23848 33232 23860
rect 32907 23820 33232 23848
rect 32907 23817 32919 23820
rect 32861 23811 32919 23817
rect 33226 23808 33232 23820
rect 33284 23808 33290 23860
rect 36814 23848 36820 23860
rect 36775 23820 36820 23848
rect 36814 23808 36820 23820
rect 36872 23808 36878 23860
rect 27890 23740 27896 23792
rect 27948 23740 27954 23792
rect 30466 23740 30472 23792
rect 30524 23740 30530 23792
rect 35434 23780 35440 23792
rect 35084 23752 35440 23780
rect 22830 23712 22836 23724
rect 22066 23684 22836 23712
rect 22830 23672 22836 23684
rect 22888 23672 22894 23724
rect 24489 23715 24547 23721
rect 24489 23681 24501 23715
rect 24535 23712 24547 23715
rect 29733 23715 29791 23721
rect 24535 23684 26096 23712
rect 24535 23681 24547 23684
rect 24489 23675 24547 23681
rect 26068 23656 26096 23684
rect 29733 23681 29745 23715
rect 29779 23712 29791 23715
rect 32490 23712 32496 23724
rect 29779 23684 30236 23712
rect 32451 23684 32496 23712
rect 29779 23681 29791 23684
rect 29733 23675 29791 23681
rect 13998 23644 14004 23656
rect 12084 23616 14004 23644
rect 11977 23607 12035 23613
rect 9582 23536 9588 23588
rect 9640 23576 9646 23588
rect 11992 23576 12020 23607
rect 13998 23604 14004 23616
rect 14056 23604 14062 23656
rect 15657 23647 15715 23653
rect 15657 23613 15669 23647
rect 15703 23613 15715 23647
rect 15657 23607 15715 23613
rect 17497 23647 17555 23653
rect 17497 23613 17509 23647
rect 17543 23644 17555 23647
rect 19702 23644 19708 23656
rect 17543 23616 19708 23644
rect 17543 23613 17555 23616
rect 17497 23607 17555 23613
rect 12342 23576 12348 23588
rect 9640 23548 12348 23576
rect 9640 23536 9646 23548
rect 12342 23536 12348 23548
rect 12400 23536 12406 23588
rect 9217 23511 9275 23517
rect 9217 23477 9229 23511
rect 9263 23508 9275 23511
rect 9306 23508 9312 23520
rect 9263 23480 9312 23508
rect 9263 23477 9275 23480
rect 9217 23471 9275 23477
rect 9306 23468 9312 23480
rect 9364 23468 9370 23520
rect 10413 23511 10471 23517
rect 10413 23477 10425 23511
rect 10459 23508 10471 23511
rect 10594 23508 10600 23520
rect 10459 23480 10600 23508
rect 10459 23477 10471 23480
rect 10413 23471 10471 23477
rect 10594 23468 10600 23480
rect 10652 23468 10658 23520
rect 12526 23508 12532 23520
rect 12487 23480 12532 23508
rect 12526 23468 12532 23480
rect 12584 23468 12590 23520
rect 15672 23508 15700 23607
rect 19702 23604 19708 23616
rect 19760 23604 19766 23656
rect 23109 23647 23167 23653
rect 23109 23613 23121 23647
rect 23155 23644 23167 23647
rect 23842 23644 23848 23656
rect 23155 23616 23848 23644
rect 23155 23613 23167 23616
rect 23109 23607 23167 23613
rect 23842 23604 23848 23616
rect 23900 23644 23906 23656
rect 24670 23644 24676 23656
rect 23900 23616 24676 23644
rect 23900 23604 23906 23616
rect 24670 23604 24676 23616
rect 24728 23604 24734 23656
rect 25682 23604 25688 23656
rect 25740 23644 25746 23656
rect 25866 23644 25872 23656
rect 25740 23616 25872 23644
rect 25740 23604 25746 23616
rect 25866 23604 25872 23616
rect 25924 23604 25930 23656
rect 26050 23644 26056 23656
rect 26011 23616 26056 23644
rect 26050 23604 26056 23616
rect 26108 23604 26114 23656
rect 27154 23644 27160 23656
rect 27115 23616 27160 23644
rect 27154 23604 27160 23616
rect 27212 23604 27218 23656
rect 27430 23644 27436 23656
rect 27391 23616 27436 23644
rect 27430 23604 27436 23616
rect 27488 23604 27494 23656
rect 30098 23644 30104 23656
rect 30059 23616 30104 23644
rect 30098 23604 30104 23616
rect 30156 23604 30162 23656
rect 30208 23644 30236 23684
rect 32490 23672 32496 23684
rect 32548 23672 32554 23724
rect 33502 23712 33508 23724
rect 33463 23684 33508 23712
rect 33502 23672 33508 23684
rect 33560 23672 33566 23724
rect 34422 23712 34428 23724
rect 34383 23684 34428 23712
rect 34422 23672 34428 23684
rect 34480 23672 34486 23724
rect 34974 23712 34980 23724
rect 34532 23684 34980 23712
rect 31938 23644 31944 23656
rect 30208 23616 31944 23644
rect 31938 23604 31944 23616
rect 31996 23604 32002 23656
rect 32398 23644 32404 23656
rect 32359 23616 32404 23644
rect 32398 23604 32404 23616
rect 32456 23604 32462 23656
rect 33594 23644 33600 23656
rect 33555 23616 33600 23644
rect 33594 23604 33600 23616
rect 33652 23604 33658 23656
rect 33873 23647 33931 23653
rect 33873 23613 33885 23647
rect 33919 23644 33931 23647
rect 34532 23644 34560 23684
rect 34974 23672 34980 23684
rect 35032 23672 35038 23724
rect 35084 23721 35112 23752
rect 35434 23740 35440 23752
rect 35492 23740 35498 23792
rect 35069 23715 35127 23721
rect 35069 23681 35081 23715
rect 35115 23681 35127 23715
rect 35069 23675 35127 23681
rect 36446 23672 36452 23724
rect 36504 23672 36510 23724
rect 35345 23647 35403 23653
rect 35345 23644 35357 23647
rect 33919 23616 34560 23644
rect 34624 23616 35357 23644
rect 33919 23613 33931 23616
rect 33873 23607 33931 23613
rect 34624 23585 34652 23616
rect 35345 23613 35357 23616
rect 35391 23613 35403 23647
rect 35345 23607 35403 23613
rect 34609 23579 34667 23585
rect 34609 23545 34621 23579
rect 34655 23545 34667 23579
rect 34609 23539 34667 23545
rect 16206 23508 16212 23520
rect 15672 23480 16212 23508
rect 16206 23468 16212 23480
rect 16264 23508 16270 23520
rect 20162 23508 20168 23520
rect 16264 23480 20168 23508
rect 16264 23468 16270 23480
rect 20162 23468 20168 23480
rect 20220 23468 20226 23520
rect 21450 23508 21456 23520
rect 21411 23480 21456 23508
rect 21450 23468 21456 23480
rect 21508 23468 21514 23520
rect 26326 23468 26332 23520
rect 26384 23508 26390 23520
rect 26513 23511 26571 23517
rect 26513 23508 26525 23511
rect 26384 23480 26525 23508
rect 26384 23468 26390 23480
rect 26513 23477 26525 23480
rect 26559 23477 26571 23511
rect 26513 23471 26571 23477
rect 31527 23511 31585 23517
rect 31527 23477 31539 23511
rect 31573 23508 31585 23511
rect 32122 23508 32128 23520
rect 31573 23480 32128 23508
rect 31573 23477 31585 23480
rect 31527 23471 31585 23477
rect 32122 23468 32128 23480
rect 32180 23508 32186 23520
rect 32306 23508 32312 23520
rect 32180 23480 32312 23508
rect 32180 23468 32186 23480
rect 32306 23468 32312 23480
rect 32364 23468 32370 23520
rect 1104 23418 37628 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 37628 23418
rect 1104 23344 37628 23366
rect 6181 23307 6239 23313
rect 6181 23273 6193 23307
rect 6227 23304 6239 23307
rect 7282 23304 7288 23316
rect 6227 23276 7288 23304
rect 6227 23273 6239 23276
rect 6181 23267 6239 23273
rect 7282 23264 7288 23276
rect 7340 23264 7346 23316
rect 7558 23264 7564 23316
rect 7616 23304 7622 23316
rect 9125 23307 9183 23313
rect 9125 23304 9137 23307
rect 7616 23276 9137 23304
rect 7616 23264 7622 23276
rect 9125 23273 9137 23276
rect 9171 23273 9183 23307
rect 9125 23267 9183 23273
rect 11330 23264 11336 23316
rect 11388 23304 11394 23316
rect 12713 23307 12771 23313
rect 12713 23304 12725 23307
rect 11388 23276 12725 23304
rect 11388 23264 11394 23276
rect 12713 23273 12725 23276
rect 12759 23273 12771 23307
rect 12713 23267 12771 23273
rect 13906 23264 13912 23316
rect 13964 23304 13970 23316
rect 14369 23307 14427 23313
rect 14369 23304 14381 23307
rect 13964 23276 14381 23304
rect 13964 23264 13970 23276
rect 14369 23273 14381 23276
rect 14415 23273 14427 23307
rect 14369 23267 14427 23273
rect 18506 23264 18512 23316
rect 18564 23304 18570 23316
rect 18601 23307 18659 23313
rect 18601 23304 18613 23307
rect 18564 23276 18613 23304
rect 18564 23264 18570 23276
rect 18601 23273 18613 23276
rect 18647 23273 18659 23307
rect 18601 23267 18659 23273
rect 19058 23264 19064 23316
rect 19116 23304 19122 23316
rect 19521 23307 19579 23313
rect 19521 23304 19533 23307
rect 19116 23276 19533 23304
rect 19116 23264 19122 23276
rect 19521 23273 19533 23276
rect 19567 23273 19579 23307
rect 19521 23267 19579 23273
rect 19610 23264 19616 23316
rect 19668 23304 19674 23316
rect 20254 23304 20260 23316
rect 19668 23276 20260 23304
rect 19668 23264 19674 23276
rect 20254 23264 20260 23276
rect 20312 23264 20318 23316
rect 20990 23264 20996 23316
rect 21048 23304 21054 23316
rect 26513 23307 26571 23313
rect 21048 23276 26464 23304
rect 21048 23264 21054 23276
rect 9766 23236 9772 23248
rect 8036 23208 9772 23236
rect 6825 23171 6883 23177
rect 6825 23137 6837 23171
rect 6871 23168 6883 23171
rect 8036 23168 8064 23208
rect 9766 23196 9772 23208
rect 9824 23196 9830 23248
rect 12158 23196 12164 23248
rect 12216 23236 12222 23248
rect 12253 23239 12311 23245
rect 12253 23236 12265 23239
rect 12216 23208 12265 23236
rect 12216 23196 12222 23208
rect 12253 23205 12265 23208
rect 12299 23205 12311 23239
rect 12253 23199 12311 23205
rect 12434 23196 12440 23248
rect 12492 23236 12498 23248
rect 13078 23236 13084 23248
rect 12492 23208 13084 23236
rect 12492 23196 12498 23208
rect 13078 23196 13084 23208
rect 13136 23196 13142 23248
rect 26436 23236 26464 23276
rect 26513 23273 26525 23307
rect 26559 23304 26571 23307
rect 27430 23304 27436 23316
rect 26559 23276 27436 23304
rect 26559 23273 26571 23276
rect 26513 23267 26571 23273
rect 27430 23264 27436 23276
rect 27488 23264 27494 23316
rect 27801 23307 27859 23313
rect 27801 23273 27813 23307
rect 27847 23304 27859 23307
rect 27890 23304 27896 23316
rect 27847 23276 27896 23304
rect 27847 23273 27859 23276
rect 27801 23267 27859 23273
rect 27890 23264 27896 23276
rect 27948 23264 27954 23316
rect 28997 23307 29055 23313
rect 28997 23273 29009 23307
rect 29043 23304 29055 23307
rect 29086 23304 29092 23316
rect 29043 23276 29092 23304
rect 29043 23273 29055 23276
rect 28997 23267 29055 23273
rect 29086 23264 29092 23276
rect 29144 23264 29150 23316
rect 30466 23304 30472 23316
rect 30427 23276 30472 23304
rect 30466 23264 30472 23276
rect 30524 23264 30530 23316
rect 31665 23307 31723 23313
rect 31665 23273 31677 23307
rect 31711 23304 31723 23307
rect 31938 23304 31944 23316
rect 31711 23276 31944 23304
rect 31711 23273 31723 23276
rect 31665 23267 31723 23273
rect 31938 23264 31944 23276
rect 31996 23264 32002 23316
rect 32766 23264 32772 23316
rect 32824 23304 32830 23316
rect 33413 23307 33471 23313
rect 33413 23304 33425 23307
rect 32824 23276 33425 23304
rect 32824 23264 32830 23276
rect 33413 23273 33425 23276
rect 33459 23273 33471 23307
rect 33413 23267 33471 23273
rect 33502 23264 33508 23316
rect 33560 23304 33566 23316
rect 33597 23307 33655 23313
rect 33597 23304 33609 23307
rect 33560 23276 33609 23304
rect 33560 23264 33566 23276
rect 33597 23273 33609 23276
rect 33643 23273 33655 23307
rect 33597 23267 33655 23273
rect 34698 23264 34704 23316
rect 34756 23304 34762 23316
rect 35161 23307 35219 23313
rect 35161 23304 35173 23307
rect 34756 23276 35173 23304
rect 34756 23264 34762 23276
rect 35161 23273 35173 23276
rect 35207 23273 35219 23307
rect 35161 23267 35219 23273
rect 26436 23208 31754 23236
rect 6871 23140 8064 23168
rect 6871 23137 6883 23140
rect 6825 23131 6883 23137
rect 8110 23128 8116 23180
rect 8168 23168 8174 23180
rect 8389 23171 8447 23177
rect 8389 23168 8401 23171
rect 8168 23140 8401 23168
rect 8168 23128 8174 23140
rect 8389 23137 8401 23140
rect 8435 23137 8447 23171
rect 8389 23131 8447 23137
rect 9582 23128 9588 23180
rect 9640 23168 9646 23180
rect 9677 23171 9735 23177
rect 9677 23168 9689 23171
rect 9640 23140 9689 23168
rect 9640 23128 9646 23140
rect 9677 23137 9689 23140
rect 9723 23137 9735 23171
rect 9677 23131 9735 23137
rect 10505 23171 10563 23177
rect 10505 23137 10517 23171
rect 10551 23168 10563 23171
rect 11514 23168 11520 23180
rect 10551 23140 11520 23168
rect 10551 23137 10563 23140
rect 10505 23131 10563 23137
rect 11514 23128 11520 23140
rect 11572 23128 11578 23180
rect 11790 23128 11796 23180
rect 11848 23168 11854 23180
rect 13170 23168 13176 23180
rect 11848 23140 12434 23168
rect 13131 23140 13176 23168
rect 11848 23128 11854 23140
rect 5997 23103 6055 23109
rect 5997 23069 6009 23103
rect 6043 23100 6055 23103
rect 8297 23103 8355 23109
rect 6043 23072 7696 23100
rect 6043 23069 6055 23072
rect 5997 23063 6055 23069
rect 7009 23035 7067 23041
rect 7009 23001 7021 23035
rect 7055 23032 7067 23035
rect 7558 23032 7564 23044
rect 7055 23004 7564 23032
rect 7055 23001 7067 23004
rect 7009 22995 7067 23001
rect 7558 22992 7564 23004
rect 7616 22992 7622 23044
rect 6914 22924 6920 22976
rect 6972 22964 6978 22976
rect 7377 22967 7435 22973
rect 6972 22936 7017 22964
rect 6972 22924 6978 22936
rect 7377 22933 7389 22967
rect 7423 22964 7435 22967
rect 7466 22964 7472 22976
rect 7423 22936 7472 22964
rect 7423 22933 7435 22936
rect 7377 22927 7435 22933
rect 7466 22924 7472 22936
rect 7524 22924 7530 22976
rect 7668 22964 7696 23072
rect 8297 23069 8309 23103
rect 8343 23100 8355 23103
rect 8570 23100 8576 23112
rect 8343 23072 8576 23100
rect 8343 23069 8355 23072
rect 8297 23063 8355 23069
rect 8570 23060 8576 23072
rect 8628 23100 8634 23112
rect 9493 23103 9551 23109
rect 9493 23100 9505 23103
rect 8628 23072 9505 23100
rect 8628 23060 8634 23072
rect 9493 23069 9505 23072
rect 9539 23069 9551 23103
rect 9493 23063 9551 23069
rect 10778 23032 10784 23044
rect 10739 23004 10784 23032
rect 10778 22992 10784 23004
rect 10836 22992 10842 23044
rect 12066 23032 12072 23044
rect 12006 23004 12072 23032
rect 12066 22992 12072 23004
rect 12124 22992 12130 23044
rect 12406 23032 12434 23140
rect 13170 23128 13176 23140
rect 13228 23128 13234 23180
rect 13265 23171 13323 23177
rect 13265 23137 13277 23171
rect 13311 23137 13323 23171
rect 13265 23131 13323 23137
rect 12526 23060 12532 23112
rect 12584 23100 12590 23112
rect 13081 23103 13139 23109
rect 13081 23100 13093 23103
rect 12584 23072 13093 23100
rect 12584 23060 12590 23072
rect 13081 23069 13093 23072
rect 13127 23069 13139 23103
rect 13081 23063 13139 23069
rect 12618 23032 12624 23044
rect 12406 23004 12624 23032
rect 12618 22992 12624 23004
rect 12676 23032 12682 23044
rect 13280 23032 13308 23131
rect 15470 23128 15476 23180
rect 15528 23168 15534 23180
rect 15841 23171 15899 23177
rect 15841 23168 15853 23171
rect 15528 23140 15853 23168
rect 15528 23128 15534 23140
rect 15841 23137 15853 23140
rect 15887 23137 15899 23171
rect 15841 23131 15899 23137
rect 16117 23171 16175 23177
rect 16117 23137 16129 23171
rect 16163 23168 16175 23171
rect 17586 23168 17592 23180
rect 16163 23140 17592 23168
rect 16163 23137 16175 23140
rect 16117 23131 16175 23137
rect 17586 23128 17592 23140
rect 17644 23128 17650 23180
rect 19886 23128 19892 23180
rect 19944 23168 19950 23180
rect 19981 23171 20039 23177
rect 19981 23168 19993 23171
rect 19944 23140 19993 23168
rect 19944 23128 19950 23140
rect 19981 23137 19993 23140
rect 20027 23137 20039 23171
rect 19981 23131 20039 23137
rect 16758 23100 16764 23112
rect 16719 23072 16764 23100
rect 16758 23060 16764 23072
rect 16816 23060 16822 23112
rect 17221 23103 17279 23109
rect 17221 23069 17233 23103
rect 17267 23100 17279 23103
rect 17494 23100 17500 23112
rect 17267 23072 17500 23100
rect 17267 23069 17279 23072
rect 17221 23063 17279 23069
rect 17494 23060 17500 23072
rect 17552 23060 17558 23112
rect 17954 23060 17960 23112
rect 18012 23100 18018 23112
rect 18509 23103 18567 23109
rect 18509 23100 18521 23103
rect 18012 23072 18521 23100
rect 18012 23060 18018 23072
rect 18509 23069 18521 23072
rect 18555 23100 18567 23103
rect 19242 23100 19248 23112
rect 18555 23072 19248 23100
rect 18555 23069 18567 23072
rect 18509 23063 18567 23069
rect 19242 23060 19248 23072
rect 19300 23060 19306 23112
rect 19996 23100 20024 23131
rect 20162 23128 20168 23180
rect 20220 23168 20226 23180
rect 20990 23168 20996 23180
rect 20220 23140 20996 23168
rect 20220 23128 20226 23140
rect 20990 23128 20996 23140
rect 21048 23128 21054 23180
rect 21637 23171 21695 23177
rect 21637 23137 21649 23171
rect 21683 23168 21695 23171
rect 21818 23168 21824 23180
rect 21683 23140 21824 23168
rect 21683 23137 21695 23140
rect 21637 23131 21695 23137
rect 21818 23128 21824 23140
rect 21876 23128 21882 23180
rect 22281 23171 22339 23177
rect 22281 23137 22293 23171
rect 22327 23168 22339 23171
rect 22646 23168 22652 23180
rect 22327 23140 22652 23168
rect 22327 23137 22339 23140
rect 22281 23131 22339 23137
rect 22646 23128 22652 23140
rect 22704 23128 22710 23180
rect 24029 23171 24087 23177
rect 24029 23137 24041 23171
rect 24075 23168 24087 23171
rect 25590 23168 25596 23180
rect 24075 23140 25452 23168
rect 25551 23140 25596 23168
rect 24075 23137 24087 23140
rect 24029 23131 24087 23137
rect 21450 23100 21456 23112
rect 19996 23072 21456 23100
rect 21450 23060 21456 23072
rect 21508 23060 21514 23112
rect 25424 23109 25452 23140
rect 25590 23128 25596 23140
rect 25648 23128 25654 23180
rect 25409 23103 25467 23109
rect 25409 23069 25421 23103
rect 25455 23100 25467 23103
rect 26050 23100 26056 23112
rect 25455 23072 26056 23100
rect 25455 23069 25467 23072
rect 25409 23063 25467 23069
rect 26050 23060 26056 23072
rect 26108 23060 26114 23112
rect 26326 23100 26332 23112
rect 26287 23072 26332 23100
rect 26326 23060 26332 23072
rect 26384 23060 26390 23112
rect 27706 23100 27712 23112
rect 27667 23072 27712 23100
rect 27706 23060 27712 23072
rect 27764 23060 27770 23112
rect 28828 23109 28856 23208
rect 31726 23168 31754 23208
rect 32490 23168 32496 23180
rect 29840 23140 30788 23168
rect 31726 23140 32496 23168
rect 28721 23103 28779 23109
rect 28721 23100 28733 23103
rect 27816 23072 28733 23100
rect 21361 23035 21419 23041
rect 12676 23004 13308 23032
rect 15410 23004 15700 23032
rect 12676 22992 12682 23004
rect 7837 22967 7895 22973
rect 7837 22964 7849 22967
rect 7668 22936 7849 22964
rect 7837 22933 7849 22936
rect 7883 22933 7895 22967
rect 7837 22927 7895 22933
rect 8205 22967 8263 22973
rect 8205 22933 8217 22967
rect 8251 22964 8263 22967
rect 8754 22964 8760 22976
rect 8251 22936 8760 22964
rect 8251 22933 8263 22936
rect 8205 22927 8263 22933
rect 8754 22924 8760 22936
rect 8812 22924 8818 22976
rect 9214 22924 9220 22976
rect 9272 22964 9278 22976
rect 9585 22967 9643 22973
rect 9585 22964 9597 22967
rect 9272 22936 9597 22964
rect 9272 22924 9278 22936
rect 9585 22933 9597 22936
rect 9631 22964 9643 22967
rect 13906 22964 13912 22976
rect 9631 22936 13912 22964
rect 9631 22933 9643 22936
rect 9585 22927 9643 22933
rect 13906 22924 13912 22936
rect 13964 22924 13970 22976
rect 15672 22964 15700 23004
rect 21361 23001 21373 23035
rect 21407 23032 21419 23035
rect 22554 23032 22560 23044
rect 21407 23004 22094 23032
rect 22515 23004 22560 23032
rect 21407 23001 21419 23004
rect 21361 22995 21419 23001
rect 16669 22967 16727 22973
rect 16669 22964 16681 22967
rect 15672 22936 16681 22964
rect 16669 22933 16681 22936
rect 16715 22933 16727 22967
rect 17310 22964 17316 22976
rect 17271 22936 17316 22964
rect 16669 22927 16727 22933
rect 17310 22924 17316 22936
rect 17368 22924 17374 22976
rect 19886 22964 19892 22976
rect 19847 22936 19892 22964
rect 19886 22924 19892 22936
rect 19944 22924 19950 22976
rect 20898 22924 20904 22976
rect 20956 22964 20962 22976
rect 20993 22967 21051 22973
rect 20993 22964 21005 22967
rect 20956 22936 21005 22964
rect 20956 22924 20962 22936
rect 20993 22933 21005 22936
rect 21039 22933 21051 22967
rect 22066 22964 22094 23004
rect 22554 22992 22560 23004
rect 22612 22992 22618 23044
rect 23566 22992 23572 23044
rect 23624 22992 23630 23044
rect 27816 23032 27844 23072
rect 28721 23069 28733 23072
rect 28767 23069 28779 23103
rect 28721 23063 28779 23069
rect 28813 23103 28871 23109
rect 28813 23069 28825 23103
rect 28859 23069 28871 23103
rect 29730 23100 29736 23112
rect 29691 23072 29736 23100
rect 28813 23063 28871 23069
rect 28442 23032 28448 23044
rect 24964 23004 27844 23032
rect 28403 23004 28448 23032
rect 24964 22964 24992 23004
rect 28442 22992 28448 23004
rect 28500 22992 28506 23044
rect 28736 23032 28764 23063
rect 29730 23060 29736 23072
rect 29788 23060 29794 23112
rect 29840 23032 29868 23140
rect 29917 23103 29975 23109
rect 29917 23069 29929 23103
rect 29963 23069 29975 23103
rect 29917 23063 29975 23069
rect 30377 23103 30435 23109
rect 30377 23069 30389 23103
rect 30423 23100 30435 23103
rect 30558 23100 30564 23112
rect 30423 23072 30564 23100
rect 30423 23069 30435 23072
rect 30377 23063 30435 23069
rect 28736 23004 29868 23032
rect 29932 23032 29960 23063
rect 30558 23060 30564 23072
rect 30616 23060 30622 23112
rect 30650 23032 30656 23044
rect 29932 23004 30656 23032
rect 30650 22992 30656 23004
rect 30708 22992 30714 23044
rect 30760 23032 30788 23140
rect 32490 23128 32496 23140
rect 32548 23128 32554 23180
rect 35434 23128 35440 23180
rect 35492 23168 35498 23180
rect 36909 23171 36967 23177
rect 36909 23168 36921 23171
rect 35492 23140 36921 23168
rect 35492 23128 35498 23140
rect 36909 23137 36921 23140
rect 36955 23137 36967 23171
rect 36909 23131 36967 23137
rect 33594 23100 33600 23112
rect 33555 23072 33600 23100
rect 33594 23060 33600 23072
rect 33652 23060 33658 23112
rect 33778 23060 33784 23112
rect 33836 23100 33842 23112
rect 33836 23072 33881 23100
rect 33836 23060 33842 23072
rect 32214 23032 32220 23044
rect 30760 23004 32220 23032
rect 32214 22992 32220 23004
rect 32272 22992 32278 23044
rect 32950 23032 32956 23044
rect 32911 23004 32956 23032
rect 32950 22992 32956 23004
rect 33008 22992 33014 23044
rect 35342 22992 35348 23044
rect 35400 23032 35406 23044
rect 36633 23035 36691 23041
rect 35400 23004 35466 23032
rect 35400 22992 35406 23004
rect 36633 23001 36645 23035
rect 36679 23001 36691 23035
rect 36633 22995 36691 23001
rect 22066 22936 24992 22964
rect 25041 22967 25099 22973
rect 20993 22927 21051 22933
rect 25041 22933 25053 22967
rect 25087 22964 25099 22967
rect 25314 22964 25320 22976
rect 25087 22936 25320 22964
rect 25087 22933 25099 22936
rect 25041 22927 25099 22933
rect 25314 22924 25320 22936
rect 25372 22924 25378 22976
rect 25501 22967 25559 22973
rect 25501 22933 25513 22967
rect 25547 22964 25559 22967
rect 25958 22964 25964 22976
rect 25547 22936 25964 22964
rect 25547 22933 25559 22936
rect 25501 22927 25559 22933
rect 25958 22924 25964 22936
rect 26016 22964 26022 22976
rect 27982 22964 27988 22976
rect 26016 22936 27988 22964
rect 26016 22924 26022 22936
rect 27982 22924 27988 22936
rect 28040 22924 28046 22976
rect 28626 22964 28632 22976
rect 28587 22936 28632 22964
rect 28626 22924 28632 22936
rect 28684 22924 28690 22976
rect 29822 22964 29828 22976
rect 29783 22936 29828 22964
rect 29822 22924 29828 22936
rect 29880 22924 29886 22976
rect 30558 22924 30564 22976
rect 30616 22964 30622 22976
rect 31110 22964 31116 22976
rect 30616 22936 31116 22964
rect 30616 22924 30622 22936
rect 31110 22924 31116 22936
rect 31168 22924 31174 22976
rect 35986 22924 35992 22976
rect 36044 22964 36050 22976
rect 36648 22964 36676 22995
rect 36044 22936 36676 22964
rect 36044 22924 36050 22936
rect 1104 22874 37628 22896
rect 1104 22822 4874 22874
rect 4926 22822 4938 22874
rect 4990 22822 5002 22874
rect 5054 22822 5066 22874
rect 5118 22822 5130 22874
rect 5182 22822 35594 22874
rect 35646 22822 35658 22874
rect 35710 22822 35722 22874
rect 35774 22822 35786 22874
rect 35838 22822 35850 22874
rect 35902 22822 37628 22874
rect 1104 22800 37628 22822
rect 6914 22720 6920 22772
rect 6972 22760 6978 22772
rect 8202 22760 8208 22772
rect 6972 22732 8208 22760
rect 6972 22720 6978 22732
rect 8202 22720 8208 22732
rect 8260 22760 8266 22772
rect 8389 22763 8447 22769
rect 8389 22760 8401 22763
rect 8260 22732 8401 22760
rect 8260 22720 8266 22732
rect 8389 22729 8401 22732
rect 8435 22729 8447 22763
rect 8389 22723 8447 22729
rect 9674 22720 9680 22772
rect 9732 22760 9738 22772
rect 10873 22763 10931 22769
rect 10873 22760 10885 22763
rect 9732 22732 10885 22760
rect 9732 22720 9738 22732
rect 10873 22729 10885 22732
rect 10919 22729 10931 22763
rect 10873 22723 10931 22729
rect 13262 22720 13268 22772
rect 13320 22760 13326 22772
rect 13449 22763 13507 22769
rect 13449 22760 13461 22763
rect 13320 22732 13461 22760
rect 13320 22720 13326 22732
rect 13449 22729 13461 22732
rect 13495 22729 13507 22763
rect 21910 22760 21916 22772
rect 13449 22723 13507 22729
rect 16132 22732 21916 22760
rect 6822 22692 6828 22704
rect 6656 22664 6828 22692
rect 6656 22633 6684 22664
rect 6822 22652 6828 22664
rect 6880 22652 6886 22704
rect 10042 22652 10048 22704
rect 10100 22652 10106 22704
rect 11882 22652 11888 22704
rect 11940 22692 11946 22704
rect 11977 22695 12035 22701
rect 11977 22692 11989 22695
rect 11940 22664 11989 22692
rect 11940 22652 11946 22664
rect 11977 22661 11989 22664
rect 12023 22661 12035 22695
rect 11977 22655 12035 22661
rect 12434 22652 12440 22704
rect 12492 22652 12498 22704
rect 14642 22652 14648 22704
rect 14700 22692 14706 22704
rect 14918 22692 14924 22704
rect 14700 22664 14924 22692
rect 14700 22652 14706 22664
rect 14918 22652 14924 22664
rect 14976 22652 14982 22704
rect 6641 22627 6699 22633
rect 6641 22593 6653 22627
rect 6687 22593 6699 22627
rect 6641 22587 6699 22593
rect 8018 22584 8024 22636
rect 8076 22584 8082 22636
rect 9122 22624 9128 22636
rect 9083 22596 9128 22624
rect 9122 22584 9128 22596
rect 9180 22584 9186 22636
rect 11698 22624 11704 22636
rect 11659 22596 11704 22624
rect 11698 22584 11704 22596
rect 11756 22584 11762 22636
rect 13906 22624 13912 22636
rect 13867 22596 13912 22624
rect 13906 22584 13912 22596
rect 13964 22584 13970 22636
rect 16132 22633 16160 22732
rect 21910 22720 21916 22732
rect 21968 22720 21974 22772
rect 25314 22760 25320 22772
rect 25275 22732 25320 22760
rect 25314 22720 25320 22732
rect 25372 22720 25378 22772
rect 26329 22763 26387 22769
rect 26329 22729 26341 22763
rect 26375 22760 26387 22763
rect 26375 22732 27476 22760
rect 26375 22729 26387 22732
rect 26329 22723 26387 22729
rect 17310 22652 17316 22704
rect 17368 22652 17374 22704
rect 23658 22652 23664 22704
rect 23716 22652 23722 22704
rect 27448 22701 27476 22732
rect 28074 22720 28080 22772
rect 28132 22760 28138 22772
rect 28905 22763 28963 22769
rect 28905 22760 28917 22763
rect 28132 22732 28917 22760
rect 28132 22720 28138 22732
rect 28905 22729 28917 22732
rect 28951 22729 28963 22763
rect 33134 22760 33140 22772
rect 28905 22723 28963 22729
rect 30576 22732 33140 22760
rect 27433 22695 27491 22701
rect 27433 22661 27445 22695
rect 27479 22661 27491 22695
rect 27433 22655 27491 22661
rect 27890 22652 27896 22704
rect 27948 22652 27954 22704
rect 16117 22627 16175 22633
rect 16117 22593 16129 22627
rect 16163 22593 16175 22627
rect 16117 22587 16175 22593
rect 18598 22584 18604 22636
rect 18656 22624 18662 22636
rect 18656 22596 18701 22624
rect 18656 22584 18662 22596
rect 19242 22584 19248 22636
rect 19300 22624 19306 22636
rect 19337 22627 19395 22633
rect 19337 22624 19349 22627
rect 19300 22596 19349 22624
rect 19300 22584 19306 22596
rect 19337 22593 19349 22596
rect 19383 22593 19395 22627
rect 20530 22624 20536 22636
rect 20491 22596 20536 22624
rect 19337 22587 19395 22593
rect 20530 22584 20536 22596
rect 20588 22584 20594 22636
rect 21174 22584 21180 22636
rect 21232 22624 21238 22636
rect 22005 22627 22063 22633
rect 22005 22624 22017 22627
rect 21232 22596 22017 22624
rect 21232 22584 21238 22596
rect 22005 22593 22017 22596
rect 22051 22593 22063 22627
rect 22738 22624 22744 22636
rect 22699 22596 22744 22624
rect 22005 22587 22063 22593
rect 22738 22584 22744 22596
rect 22796 22584 22802 22636
rect 24670 22584 24676 22636
rect 24728 22624 24734 22636
rect 26142 22624 26148 22636
rect 24728 22596 25544 22624
rect 26103 22596 26148 22624
rect 24728 22584 24734 22596
rect 6914 22516 6920 22568
rect 6972 22556 6978 22568
rect 9398 22556 9404 22568
rect 6972 22528 7017 22556
rect 9359 22528 9404 22556
rect 6972 22516 6978 22528
rect 9398 22516 9404 22528
rect 9456 22516 9462 22568
rect 18325 22559 18383 22565
rect 18325 22556 18337 22559
rect 16316 22528 18337 22556
rect 13998 22448 14004 22500
rect 14056 22488 14062 22500
rect 15197 22491 15255 22497
rect 14056 22460 15148 22488
rect 14056 22448 14062 22460
rect 14090 22420 14096 22432
rect 14051 22392 14096 22420
rect 14090 22380 14096 22392
rect 14148 22380 14154 22432
rect 15120 22420 15148 22460
rect 15197 22457 15209 22491
rect 15243 22488 15255 22491
rect 15562 22488 15568 22500
rect 15243 22460 15568 22488
rect 15243 22457 15255 22460
rect 15197 22451 15255 22457
rect 15562 22448 15568 22460
rect 15620 22448 15626 22500
rect 16316 22497 16344 22528
rect 18325 22525 18337 22528
rect 18371 22525 18383 22559
rect 18325 22519 18383 22525
rect 19886 22516 19892 22568
rect 19944 22556 19950 22568
rect 20625 22559 20683 22565
rect 20625 22556 20637 22559
rect 19944 22528 20637 22556
rect 19944 22516 19950 22528
rect 20625 22525 20637 22528
rect 20671 22525 20683 22559
rect 20625 22519 20683 22525
rect 20717 22559 20775 22565
rect 20717 22525 20729 22559
rect 20763 22525 20775 22559
rect 23014 22556 23020 22568
rect 22975 22528 23020 22556
rect 20717 22519 20775 22525
rect 16301 22491 16359 22497
rect 16301 22457 16313 22491
rect 16347 22457 16359 22491
rect 16301 22451 16359 22457
rect 20254 22448 20260 22500
rect 20312 22488 20318 22500
rect 20732 22488 20760 22519
rect 23014 22516 23020 22528
rect 23072 22516 23078 22568
rect 24489 22559 24547 22565
rect 24489 22525 24501 22559
rect 24535 22556 24547 22559
rect 25406 22556 25412 22568
rect 24535 22528 25412 22556
rect 24535 22525 24547 22528
rect 24489 22519 24547 22525
rect 25406 22516 25412 22528
rect 25464 22516 25470 22568
rect 25516 22565 25544 22596
rect 26142 22584 26148 22596
rect 26200 22584 26206 22636
rect 30576 22633 30604 22732
rect 33134 22720 33140 22732
rect 33192 22720 33198 22772
rect 35897 22763 35955 22769
rect 35897 22729 35909 22763
rect 35943 22760 35955 22763
rect 35986 22760 35992 22772
rect 35943 22732 35992 22760
rect 35943 22729 35955 22732
rect 35897 22723 35955 22729
rect 35986 22720 35992 22732
rect 36044 22720 36050 22772
rect 36446 22760 36452 22772
rect 36407 22732 36452 22760
rect 36446 22720 36452 22732
rect 36504 22720 36510 22772
rect 30650 22652 30656 22704
rect 30708 22692 30714 22704
rect 30708 22664 30753 22692
rect 30708 22652 30714 22664
rect 31754 22652 31760 22704
rect 31812 22692 31818 22704
rect 32677 22695 32735 22701
rect 32677 22692 32689 22695
rect 31812 22664 32689 22692
rect 31812 22652 31818 22664
rect 32677 22661 32689 22664
rect 32723 22661 32735 22695
rect 32677 22655 32735 22661
rect 32766 22652 32772 22704
rect 32824 22701 32830 22704
rect 32824 22695 32853 22701
rect 32841 22661 32853 22695
rect 32824 22655 32853 22661
rect 32824 22652 32830 22655
rect 32950 22652 32956 22704
rect 33008 22692 33014 22704
rect 33505 22695 33563 22701
rect 33505 22692 33517 22695
rect 33008 22664 33517 22692
rect 33008 22652 33014 22664
rect 33505 22661 33517 22664
rect 33551 22661 33563 22695
rect 33505 22655 33563 22661
rect 35253 22695 35311 22701
rect 35253 22661 35265 22695
rect 35299 22692 35311 22695
rect 36078 22692 36084 22704
rect 35299 22664 36084 22692
rect 35299 22661 35311 22664
rect 35253 22655 35311 22661
rect 36078 22652 36084 22664
rect 36136 22652 36142 22704
rect 29917 22627 29975 22633
rect 29917 22593 29929 22627
rect 29963 22624 29975 22627
rect 30561 22627 30619 22633
rect 30561 22624 30573 22627
rect 29963 22596 30573 22624
rect 29963 22593 29975 22596
rect 29917 22587 29975 22593
rect 30561 22593 30573 22596
rect 30607 22593 30619 22627
rect 30742 22624 30748 22636
rect 30703 22596 30748 22624
rect 30561 22587 30619 22593
rect 30742 22584 30748 22596
rect 30800 22584 30806 22636
rect 32493 22627 32551 22633
rect 32493 22593 32505 22627
rect 32539 22593 32551 22627
rect 32493 22587 32551 22593
rect 32585 22627 32643 22633
rect 32585 22593 32597 22627
rect 32631 22624 32643 22627
rect 33686 22624 33692 22636
rect 32631 22596 33692 22624
rect 32631 22593 32643 22596
rect 32585 22587 32643 22593
rect 25501 22559 25559 22565
rect 25501 22525 25513 22559
rect 25547 22525 25559 22559
rect 27154 22556 27160 22568
rect 27115 22528 27160 22556
rect 25501 22519 25559 22525
rect 27154 22516 27160 22528
rect 27212 22516 27218 22568
rect 30101 22559 30159 22565
rect 30101 22525 30113 22559
rect 30147 22556 30159 22559
rect 30760 22556 30788 22584
rect 30147 22528 30788 22556
rect 30147 22525 30159 22528
rect 30101 22519 30159 22525
rect 20312 22460 20760 22488
rect 20312 22448 20318 22460
rect 30374 22448 30380 22500
rect 30432 22488 30438 22500
rect 32508 22488 32536 22587
rect 33686 22584 33692 22596
rect 33744 22584 33750 22636
rect 35713 22627 35771 22633
rect 35713 22624 35725 22627
rect 35268 22596 35725 22624
rect 35268 22568 35296 22596
rect 35713 22593 35725 22596
rect 35759 22593 35771 22627
rect 36538 22624 36544 22636
rect 36499 22596 36544 22624
rect 35713 22587 35771 22593
rect 36538 22584 36544 22596
rect 36596 22584 36602 22636
rect 32953 22559 33011 22565
rect 32953 22525 32965 22559
rect 32999 22556 33011 22559
rect 33134 22556 33140 22568
rect 32999 22528 33140 22556
rect 32999 22525 33011 22528
rect 32953 22519 33011 22525
rect 33134 22516 33140 22528
rect 33192 22516 33198 22568
rect 35250 22516 35256 22568
rect 35308 22516 35314 22568
rect 33962 22488 33968 22500
rect 30432 22460 31754 22488
rect 32508 22460 33968 22488
rect 30432 22448 30438 22460
rect 16853 22423 16911 22429
rect 16853 22420 16865 22423
rect 15120 22392 16865 22420
rect 16853 22389 16865 22392
rect 16899 22389 16911 22423
rect 16853 22383 16911 22389
rect 17586 22380 17592 22432
rect 17644 22420 17650 22432
rect 18598 22420 18604 22432
rect 17644 22392 18604 22420
rect 17644 22380 17650 22392
rect 18598 22380 18604 22392
rect 18656 22380 18662 22432
rect 19242 22420 19248 22432
rect 19203 22392 19248 22420
rect 19242 22380 19248 22392
rect 19300 22380 19306 22432
rect 20162 22420 20168 22432
rect 20123 22392 20168 22420
rect 20162 22380 20168 22392
rect 20220 22380 20226 22432
rect 22094 22380 22100 22432
rect 22152 22420 22158 22432
rect 24946 22420 24952 22432
rect 22152 22392 22197 22420
rect 24907 22392 24952 22420
rect 22152 22380 22158 22392
rect 24946 22380 24952 22392
rect 25004 22380 25010 22432
rect 29730 22420 29736 22432
rect 29691 22392 29736 22420
rect 29730 22380 29736 22392
rect 29788 22380 29794 22432
rect 31726 22420 31754 22460
rect 33962 22448 33968 22460
rect 34020 22448 34026 22500
rect 32309 22423 32367 22429
rect 32309 22420 32321 22423
rect 31726 22392 32321 22420
rect 32309 22389 32321 22392
rect 32355 22389 32367 22423
rect 32309 22383 32367 22389
rect 1104 22330 37628 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 37628 22330
rect 1104 22256 37628 22278
rect 6914 22176 6920 22228
rect 6972 22216 6978 22228
rect 7285 22219 7343 22225
rect 7285 22216 7297 22219
rect 6972 22188 7297 22216
rect 6972 22176 6978 22188
rect 7285 22185 7297 22188
rect 7331 22185 7343 22219
rect 7285 22179 7343 22185
rect 9398 22176 9404 22228
rect 9456 22216 9462 22228
rect 9493 22219 9551 22225
rect 9493 22216 9505 22219
rect 9456 22188 9505 22216
rect 9456 22176 9462 22188
rect 9493 22185 9505 22188
rect 9539 22185 9551 22219
rect 10778 22216 10784 22228
rect 10739 22188 10784 22216
rect 9493 22179 9551 22185
rect 10778 22176 10784 22188
rect 10836 22176 10842 22228
rect 14090 22176 14096 22228
rect 14148 22216 14154 22228
rect 14534 22219 14592 22225
rect 14534 22216 14546 22219
rect 14148 22188 14546 22216
rect 14148 22176 14154 22188
rect 14534 22185 14546 22188
rect 14580 22185 14592 22219
rect 14534 22179 14592 22185
rect 17678 22176 17684 22228
rect 17736 22216 17742 22228
rect 20254 22216 20260 22228
rect 17736 22188 20260 22216
rect 17736 22176 17742 22188
rect 20254 22176 20260 22188
rect 20312 22176 20318 22228
rect 31938 22216 31944 22228
rect 31851 22188 31944 22216
rect 31938 22176 31944 22188
rect 31996 22216 32002 22228
rect 32582 22216 32588 22228
rect 31996 22188 32588 22216
rect 31996 22176 32002 22188
rect 32582 22176 32588 22188
rect 32640 22176 32646 22228
rect 33502 22176 33508 22228
rect 33560 22216 33566 22228
rect 34422 22216 34428 22228
rect 33560 22188 34428 22216
rect 33560 22176 33566 22188
rect 34422 22176 34428 22188
rect 34480 22176 34486 22228
rect 11698 22108 11704 22160
rect 11756 22148 11762 22160
rect 11756 22120 13676 22148
rect 11756 22108 11762 22120
rect 8018 22080 8024 22092
rect 7979 22052 8024 22080
rect 8018 22040 8024 22052
rect 8076 22040 8082 22092
rect 8294 22080 8300 22092
rect 8128 22052 8300 22080
rect 7466 22012 7472 22024
rect 7427 21984 7472 22012
rect 7466 21972 7472 21984
rect 7524 21972 7530 22024
rect 8128 22021 8156 22052
rect 8294 22040 8300 22052
rect 8352 22080 8358 22092
rect 10042 22080 10048 22092
rect 8352 22052 9536 22080
rect 10003 22052 10048 22080
rect 8352 22040 8358 22052
rect 9508 22024 9536 22052
rect 10042 22040 10048 22052
rect 10100 22040 10106 22092
rect 11977 22083 12035 22089
rect 11977 22049 11989 22083
rect 12023 22080 12035 22083
rect 12434 22080 12440 22092
rect 12023 22052 12440 22080
rect 12023 22049 12035 22052
rect 11977 22043 12035 22049
rect 12434 22040 12440 22052
rect 12492 22040 12498 22092
rect 13078 22080 13084 22092
rect 13039 22052 13084 22080
rect 13078 22040 13084 22052
rect 13136 22040 13142 22092
rect 13648 22080 13676 22120
rect 15562 22108 15568 22160
rect 15620 22148 15626 22160
rect 18966 22148 18972 22160
rect 15620 22120 18972 22148
rect 15620 22108 15626 22120
rect 13648 22052 13860 22080
rect 8113 22015 8171 22021
rect 8113 21981 8125 22015
rect 8159 21981 8171 22015
rect 9306 22012 9312 22024
rect 9267 21984 9312 22012
rect 8113 21975 8171 21981
rect 9306 21972 9312 21984
rect 9364 21972 9370 22024
rect 9490 21972 9496 22024
rect 9548 22012 9554 22024
rect 9953 22015 10011 22021
rect 9953 22012 9965 22015
rect 9548 21984 9965 22012
rect 9548 21972 9554 21984
rect 9953 21981 9965 21984
rect 9999 21981 10011 22015
rect 10594 22012 10600 22024
rect 10555 21984 10600 22012
rect 9953 21975 10011 21981
rect 10594 21972 10600 21984
rect 10652 21972 10658 22024
rect 12069 22015 12127 22021
rect 12069 21981 12081 22015
rect 12115 22012 12127 22015
rect 12158 22012 12164 22024
rect 12115 21984 12164 22012
rect 12115 21981 12127 21984
rect 12069 21975 12127 21981
rect 12158 21972 12164 21984
rect 12216 21972 12222 22024
rect 12897 22015 12955 22021
rect 12897 21981 12909 22015
rect 12943 22012 12955 22015
rect 13170 22012 13176 22024
rect 12943 21984 13176 22012
rect 12943 21981 12955 21984
rect 12897 21975 12955 21981
rect 13170 21972 13176 21984
rect 13228 21972 13234 22024
rect 13832 22012 13860 22052
rect 14918 22040 14924 22092
rect 14976 22080 14982 22092
rect 17589 22083 17647 22089
rect 14976 22052 16574 22080
rect 14976 22040 14982 22052
rect 14090 22012 14096 22024
rect 13832 21984 14096 22012
rect 14090 21972 14096 21984
rect 14148 22012 14154 22024
rect 14277 22015 14335 22021
rect 14277 22012 14289 22015
rect 14148 21984 14289 22012
rect 14148 21972 14154 21984
rect 14277 21981 14289 21984
rect 14323 21981 14335 22015
rect 14277 21975 14335 21981
rect 15010 21904 15016 21956
rect 15068 21904 15074 21956
rect 16546 21944 16574 22052
rect 17589 22049 17601 22083
rect 17635 22080 17647 22083
rect 17678 22080 17684 22092
rect 17635 22052 17684 22080
rect 17635 22049 17647 22052
rect 17589 22043 17647 22049
rect 17678 22040 17684 22052
rect 17736 22040 17742 22092
rect 18340 22089 18368 22120
rect 18966 22108 18972 22120
rect 19024 22108 19030 22160
rect 19886 22148 19892 22160
rect 19306 22120 19892 22148
rect 18325 22083 18383 22089
rect 18325 22049 18337 22083
rect 18371 22080 18383 22083
rect 18371 22052 18405 22080
rect 18371 22049 18383 22052
rect 18325 22043 18383 22049
rect 16761 22015 16819 22021
rect 16761 21981 16773 22015
rect 16807 22012 16819 22015
rect 17494 22012 17500 22024
rect 16807 21984 17500 22012
rect 16807 21981 16819 21984
rect 16761 21975 16819 21981
rect 17494 21972 17500 21984
rect 17552 21972 17558 22024
rect 18230 21972 18236 22024
rect 18288 22012 18294 22024
rect 18417 22015 18475 22021
rect 18417 22012 18429 22015
rect 18288 21984 18429 22012
rect 18288 21972 18294 21984
rect 18417 21981 18429 21984
rect 18463 22012 18475 22015
rect 19306 22012 19334 22120
rect 19886 22108 19892 22120
rect 19944 22108 19950 22160
rect 28442 22108 28448 22160
rect 28500 22148 28506 22160
rect 33594 22148 33600 22160
rect 28500 22120 33600 22148
rect 28500 22108 28506 22120
rect 19794 22040 19800 22092
rect 19852 22080 19858 22092
rect 20349 22083 20407 22089
rect 20349 22080 20361 22083
rect 19852 22052 20361 22080
rect 19852 22040 19858 22052
rect 20349 22049 20361 22052
rect 20395 22049 20407 22083
rect 20349 22043 20407 22049
rect 23293 22083 23351 22089
rect 23293 22049 23305 22083
rect 23339 22080 23351 22083
rect 23566 22080 23572 22092
rect 23339 22052 23572 22080
rect 23339 22049 23351 22052
rect 23293 22043 23351 22049
rect 23566 22040 23572 22052
rect 23624 22040 23630 22092
rect 24946 22080 24952 22092
rect 24044 22052 24952 22080
rect 18463 21984 19334 22012
rect 19705 22015 19763 22021
rect 18463 21981 18475 21984
rect 18417 21975 18475 21981
rect 19705 21981 19717 22015
rect 19751 22012 19763 22015
rect 20162 22012 20168 22024
rect 19751 21984 20168 22012
rect 19751 21981 19763 21984
rect 19705 21975 19763 21981
rect 20162 21972 20168 21984
rect 20220 21972 20226 22024
rect 22094 22012 22100 22024
rect 21758 21984 22100 22012
rect 22094 21972 22100 21984
rect 22152 21972 22158 22024
rect 24044 22021 24072 22052
rect 24946 22040 24952 22052
rect 25004 22040 25010 22092
rect 25682 22080 25688 22092
rect 25643 22052 25688 22080
rect 25682 22040 25688 22052
rect 25740 22040 25746 22092
rect 27617 22083 27675 22089
rect 27617 22049 27629 22083
rect 27663 22080 27675 22083
rect 27890 22080 27896 22092
rect 27663 22052 27896 22080
rect 27663 22049 27675 22052
rect 27617 22043 27675 22049
rect 27890 22040 27896 22052
rect 27948 22040 27954 22092
rect 28718 22080 28724 22092
rect 28679 22052 28724 22080
rect 28718 22040 28724 22052
rect 28776 22040 28782 22092
rect 30009 22083 30067 22089
rect 30009 22049 30021 22083
rect 30055 22049 30067 22083
rect 30282 22080 30288 22092
rect 30243 22052 30288 22080
rect 30009 22043 30067 22049
rect 23201 22015 23259 22021
rect 23201 21981 23213 22015
rect 23247 21981 23259 22015
rect 23201 21975 23259 21981
rect 24029 22015 24087 22021
rect 24029 21981 24041 22015
rect 24075 21981 24087 22015
rect 24029 21975 24087 21981
rect 17126 21944 17132 21956
rect 16546 21916 17132 21944
rect 17126 21904 17132 21916
rect 17184 21944 17190 21956
rect 17313 21947 17371 21953
rect 17313 21944 17325 21947
rect 17184 21916 17325 21944
rect 17184 21904 17190 21916
rect 17313 21913 17325 21916
rect 17359 21913 17371 21947
rect 20625 21947 20683 21953
rect 20625 21944 20637 21947
rect 17313 21907 17371 21913
rect 19904 21916 20637 21944
rect 12434 21836 12440 21888
rect 12492 21876 12498 21888
rect 12529 21879 12587 21885
rect 12529 21876 12541 21879
rect 12492 21848 12541 21876
rect 12492 21836 12498 21848
rect 12529 21845 12541 21848
rect 12575 21845 12587 21879
rect 12529 21839 12587 21845
rect 12802 21836 12808 21888
rect 12860 21876 12866 21888
rect 12986 21876 12992 21888
rect 12860 21848 12992 21876
rect 12860 21836 12866 21848
rect 12986 21836 12992 21848
rect 13044 21836 13050 21888
rect 16022 21876 16028 21888
rect 15983 21848 16028 21876
rect 16022 21836 16028 21848
rect 16080 21836 16086 21888
rect 16666 21876 16672 21888
rect 16627 21848 16672 21876
rect 16666 21836 16672 21848
rect 16724 21836 16730 21888
rect 18509 21879 18567 21885
rect 18509 21845 18521 21879
rect 18555 21876 18567 21879
rect 18690 21876 18696 21888
rect 18555 21848 18696 21876
rect 18555 21845 18567 21848
rect 18509 21839 18567 21845
rect 18690 21836 18696 21848
rect 18748 21836 18754 21888
rect 18874 21876 18880 21888
rect 18835 21848 18880 21876
rect 18874 21836 18880 21848
rect 18932 21836 18938 21888
rect 19904 21885 19932 21916
rect 20625 21913 20637 21916
rect 20671 21913 20683 21947
rect 23216 21944 23244 21975
rect 24486 21972 24492 22024
rect 24544 22012 24550 22024
rect 24765 22015 24823 22021
rect 24765 22012 24777 22015
rect 24544 21984 24777 22012
rect 24544 21972 24550 21984
rect 24765 21981 24777 21984
rect 24811 21981 24823 22015
rect 25958 22012 25964 22024
rect 25919 21984 25964 22012
rect 24765 21975 24823 21981
rect 25958 21972 25964 21984
rect 26016 21972 26022 22024
rect 27065 22015 27123 22021
rect 27065 21981 27077 22015
rect 27111 22012 27123 22015
rect 27525 22015 27583 22021
rect 27525 22012 27537 22015
rect 27111 21984 27537 22012
rect 27111 21981 27123 21984
rect 27065 21975 27123 21981
rect 27525 21981 27537 21984
rect 27571 22012 27583 22015
rect 27706 22012 27712 22024
rect 27571 21984 27712 22012
rect 27571 21981 27583 21984
rect 27525 21975 27583 21981
rect 27706 21972 27712 21984
rect 27764 21972 27770 22024
rect 28813 22015 28871 22021
rect 28813 21981 28825 22015
rect 28859 22012 28871 22015
rect 29362 22012 29368 22024
rect 28859 21984 29368 22012
rect 28859 21981 28871 21984
rect 28813 21975 28871 21981
rect 29362 21972 29368 21984
rect 29420 21972 29426 22024
rect 29546 21972 29552 22024
rect 29604 22012 29610 22024
rect 29822 22012 29828 22024
rect 29604 21984 29828 22012
rect 29604 21972 29610 21984
rect 29822 21972 29828 21984
rect 29880 22012 29886 22024
rect 29917 22015 29975 22021
rect 29917 22012 29929 22015
rect 29880 21984 29929 22012
rect 29880 21972 29886 21984
rect 29917 21981 29929 21984
rect 29963 21981 29975 22015
rect 30024 22012 30052 22043
rect 30282 22040 30288 22052
rect 30340 22040 30346 22092
rect 31389 22083 31447 22089
rect 31389 22049 31401 22083
rect 31435 22080 31447 22083
rect 31754 22080 31760 22092
rect 31435 22052 31760 22080
rect 31435 22049 31447 22052
rect 31389 22043 31447 22049
rect 31754 22040 31760 22052
rect 31812 22040 31818 22092
rect 30374 22012 30380 22024
rect 30024 21984 30380 22012
rect 29917 21975 29975 21981
rect 30374 21972 30380 21984
rect 30432 21972 30438 22024
rect 31113 22015 31171 22021
rect 31113 21981 31125 22015
rect 31159 21981 31171 22015
rect 31113 21975 31171 21981
rect 31205 22015 31263 22021
rect 31205 21981 31217 22015
rect 31251 22012 31263 22015
rect 31938 22012 31944 22024
rect 31251 21984 31944 22012
rect 31251 21981 31263 21984
rect 31205 21975 31263 21981
rect 23566 21944 23572 21956
rect 23216 21916 23572 21944
rect 20625 21907 20683 21913
rect 23566 21904 23572 21916
rect 23624 21904 23630 21956
rect 25406 21904 25412 21956
rect 25464 21944 25470 21956
rect 25869 21947 25927 21953
rect 25869 21944 25881 21947
rect 25464 21916 25881 21944
rect 25464 21904 25470 21916
rect 25869 21913 25881 21916
rect 25915 21913 25927 21947
rect 31128 21944 31156 21975
rect 31938 21972 31944 21984
rect 31996 21972 32002 22024
rect 32048 22012 32076 22120
rect 33594 22108 33600 22120
rect 33652 22148 33658 22160
rect 34790 22148 34796 22160
rect 33652 22120 34796 22148
rect 33652 22108 33658 22120
rect 34790 22108 34796 22120
rect 34848 22108 34854 22160
rect 32309 22083 32367 22089
rect 32309 22049 32321 22083
rect 32355 22080 32367 22083
rect 32398 22080 32404 22092
rect 32355 22052 32404 22080
rect 32355 22049 32367 22052
rect 32309 22043 32367 22049
rect 32398 22040 32404 22052
rect 32456 22040 32462 22092
rect 33686 22040 33692 22092
rect 33744 22080 33750 22092
rect 33744 22052 33824 22080
rect 33744 22040 33750 22052
rect 32217 22015 32275 22021
rect 32217 22012 32229 22015
rect 32048 21984 32229 22012
rect 32217 21981 32229 21984
rect 32263 21981 32275 22015
rect 33594 22012 33600 22024
rect 33555 21984 33600 22012
rect 32217 21975 32275 21981
rect 33594 21972 33600 21984
rect 33652 21972 33658 22024
rect 33796 22021 33824 22052
rect 34422 22040 34428 22092
rect 34480 22080 34486 22092
rect 35253 22083 35311 22089
rect 35253 22080 35265 22083
rect 34480 22052 35265 22080
rect 34480 22040 34486 22052
rect 35253 22049 35265 22052
rect 35299 22049 35311 22083
rect 35253 22043 35311 22049
rect 35342 22040 35348 22092
rect 35400 22080 35406 22092
rect 36817 22083 36875 22089
rect 36817 22080 36829 22083
rect 35400 22052 36829 22080
rect 35400 22040 35406 22052
rect 36817 22049 36829 22052
rect 36863 22049 36875 22083
rect 36817 22043 36875 22049
rect 33781 22015 33839 22021
rect 33781 21981 33793 22015
rect 33827 21981 33839 22015
rect 33962 22012 33968 22024
rect 33923 21984 33968 22012
rect 33781 21975 33839 21981
rect 33962 21972 33968 21984
rect 34020 21972 34026 22024
rect 35069 22015 35127 22021
rect 35069 21981 35081 22015
rect 35115 21981 35127 22015
rect 35069 21975 35127 21981
rect 35989 22015 36047 22021
rect 35989 21981 36001 22015
rect 36035 22012 36047 22015
rect 36078 22012 36084 22024
rect 36035 21984 36084 22012
rect 36035 21981 36047 21984
rect 35989 21975 36047 21981
rect 32858 21944 32864 21956
rect 31128 21916 32864 21944
rect 25869 21907 25927 21913
rect 32858 21904 32864 21916
rect 32916 21904 32922 21956
rect 33134 21904 33140 21956
rect 33192 21944 33198 21956
rect 33689 21947 33747 21953
rect 33689 21944 33701 21947
rect 33192 21916 33701 21944
rect 33192 21904 33198 21916
rect 33689 21913 33701 21916
rect 33735 21944 33747 21947
rect 35084 21944 35112 21975
rect 36078 21972 36084 21984
rect 36136 22012 36142 22024
rect 36538 22012 36544 22024
rect 36136 21984 36544 22012
rect 36136 21972 36142 21984
rect 36538 21972 36544 21984
rect 36596 22012 36602 22024
rect 36725 22015 36783 22021
rect 36725 22012 36737 22015
rect 36596 21984 36737 22012
rect 36596 21972 36602 21984
rect 36725 21981 36737 21984
rect 36771 21981 36783 22015
rect 36725 21975 36783 21981
rect 33735 21916 35112 21944
rect 33735 21913 33747 21916
rect 33689 21907 33747 21913
rect 19889 21879 19947 21885
rect 19889 21845 19901 21879
rect 19935 21845 19947 21879
rect 19889 21839 19947 21845
rect 22002 21836 22008 21888
rect 22060 21876 22066 21888
rect 22097 21879 22155 21885
rect 22097 21876 22109 21879
rect 22060 21848 22109 21876
rect 22060 21836 22066 21848
rect 22097 21845 22109 21848
rect 22143 21845 22155 21879
rect 22097 21839 22155 21845
rect 23014 21836 23020 21888
rect 23072 21876 23078 21888
rect 23845 21879 23903 21885
rect 23845 21876 23857 21879
rect 23072 21848 23857 21876
rect 23072 21836 23078 21848
rect 23845 21845 23857 21848
rect 23891 21845 23903 21879
rect 24670 21876 24676 21888
rect 24631 21848 24676 21876
rect 23845 21839 23903 21845
rect 24670 21836 24676 21848
rect 24728 21836 24734 21888
rect 26142 21836 26148 21888
rect 26200 21876 26206 21888
rect 26329 21879 26387 21885
rect 26329 21876 26341 21879
rect 26200 21848 26341 21876
rect 26200 21836 26206 21848
rect 26329 21845 26341 21848
rect 26375 21845 26387 21879
rect 26970 21876 26976 21888
rect 26931 21848 26976 21876
rect 26329 21839 26387 21845
rect 26970 21836 26976 21848
rect 27028 21836 27034 21888
rect 29178 21876 29184 21888
rect 29139 21848 29184 21876
rect 29178 21836 29184 21848
rect 29236 21836 29242 21888
rect 33410 21876 33416 21888
rect 33371 21848 33416 21876
rect 33410 21836 33416 21848
rect 33468 21836 33474 21888
rect 33594 21836 33600 21888
rect 33652 21876 33658 21888
rect 34885 21879 34943 21885
rect 34885 21876 34897 21879
rect 33652 21848 34897 21876
rect 33652 21836 33658 21848
rect 34885 21845 34897 21848
rect 34931 21845 34943 21879
rect 34885 21839 34943 21845
rect 35986 21836 35992 21888
rect 36044 21876 36050 21888
rect 36081 21879 36139 21885
rect 36081 21876 36093 21879
rect 36044 21848 36093 21876
rect 36044 21836 36050 21848
rect 36081 21845 36093 21848
rect 36127 21845 36139 21879
rect 36081 21839 36139 21845
rect 1104 21786 37628 21808
rect 1104 21734 4874 21786
rect 4926 21734 4938 21786
rect 4990 21734 5002 21786
rect 5054 21734 5066 21786
rect 5118 21734 5130 21786
rect 5182 21734 35594 21786
rect 35646 21734 35658 21786
rect 35710 21734 35722 21786
rect 35774 21734 35786 21786
rect 35838 21734 35850 21786
rect 35902 21734 37628 21786
rect 1104 21712 37628 21734
rect 12066 21672 12072 21684
rect 12027 21644 12072 21672
rect 12066 21632 12072 21644
rect 12124 21632 12130 21684
rect 13906 21672 13912 21684
rect 13867 21644 13912 21672
rect 13906 21632 13912 21644
rect 13964 21632 13970 21684
rect 14737 21675 14795 21681
rect 14737 21641 14749 21675
rect 14783 21672 14795 21675
rect 15010 21672 15016 21684
rect 14783 21644 15016 21672
rect 14783 21641 14795 21644
rect 14737 21635 14795 21641
rect 15010 21632 15016 21644
rect 15068 21632 15074 21684
rect 18230 21672 18236 21684
rect 18191 21644 18236 21672
rect 18230 21632 18236 21644
rect 18288 21632 18294 21684
rect 18690 21632 18696 21684
rect 18748 21672 18754 21684
rect 20441 21675 20499 21681
rect 20441 21672 20453 21675
rect 18748 21644 20453 21672
rect 18748 21632 18754 21644
rect 20441 21641 20453 21644
rect 20487 21641 20499 21675
rect 20441 21635 20499 21641
rect 20530 21632 20536 21684
rect 20588 21672 20594 21684
rect 20901 21675 20959 21681
rect 20901 21672 20913 21675
rect 20588 21644 20913 21672
rect 20588 21632 20594 21644
rect 20901 21641 20913 21644
rect 20947 21672 20959 21675
rect 22002 21672 22008 21684
rect 20947 21644 22008 21672
rect 20947 21641 20959 21644
rect 20901 21635 20959 21641
rect 22002 21632 22008 21644
rect 22060 21672 22066 21684
rect 22465 21675 22523 21681
rect 22465 21672 22477 21675
rect 22060 21644 22477 21672
rect 22060 21632 22066 21644
rect 22465 21641 22477 21644
rect 22511 21641 22523 21675
rect 23658 21672 23664 21684
rect 23619 21644 23664 21672
rect 22465 21635 22523 21641
rect 23658 21632 23664 21644
rect 23716 21632 23722 21684
rect 25406 21632 25412 21684
rect 25464 21672 25470 21684
rect 25593 21675 25651 21681
rect 25593 21672 25605 21675
rect 25464 21644 25605 21672
rect 25464 21632 25470 21644
rect 25593 21641 25605 21644
rect 25639 21641 25651 21675
rect 25593 21635 25651 21641
rect 25685 21675 25743 21681
rect 25685 21641 25697 21675
rect 25731 21672 25743 21675
rect 27246 21672 27252 21684
rect 25731 21644 27252 21672
rect 25731 21641 25743 21644
rect 25685 21635 25743 21641
rect 27246 21632 27252 21644
rect 27304 21672 27310 21684
rect 28905 21675 28963 21681
rect 28905 21672 28917 21675
rect 27304 21644 28917 21672
rect 27304 21632 27310 21644
rect 28905 21641 28917 21644
rect 28951 21641 28963 21675
rect 29546 21672 29552 21684
rect 29507 21644 29552 21672
rect 28905 21635 28963 21641
rect 29546 21632 29552 21644
rect 29604 21632 29610 21684
rect 30282 21632 30288 21684
rect 30340 21672 30346 21684
rect 30469 21675 30527 21681
rect 30469 21672 30481 21675
rect 30340 21644 30481 21672
rect 30340 21632 30346 21644
rect 30469 21641 30481 21644
rect 30515 21641 30527 21675
rect 32858 21672 32864 21684
rect 32819 21644 32864 21672
rect 30469 21635 30527 21641
rect 32858 21632 32864 21644
rect 32916 21632 32922 21684
rect 12986 21564 12992 21616
rect 13044 21604 13050 21616
rect 13541 21607 13599 21613
rect 13541 21604 13553 21607
rect 13044 21576 13553 21604
rect 13044 21564 13050 21576
rect 13541 21573 13553 21576
rect 13587 21604 13599 21607
rect 16022 21604 16028 21616
rect 13587 21576 16028 21604
rect 13587 21573 13599 21576
rect 13541 21567 13599 21573
rect 16022 21564 16028 21576
rect 16080 21564 16086 21616
rect 17494 21564 17500 21616
rect 17552 21564 17558 21616
rect 19242 21564 19248 21616
rect 19300 21564 19306 21616
rect 19794 21564 19800 21616
rect 19852 21604 19858 21616
rect 19852 21576 20024 21604
rect 19852 21564 19858 21576
rect 7837 21539 7895 21545
rect 7837 21505 7849 21539
rect 7883 21536 7895 21539
rect 8294 21536 8300 21548
rect 7883 21508 8300 21536
rect 7883 21505 7895 21508
rect 7837 21499 7895 21505
rect 8294 21496 8300 21508
rect 8352 21496 8358 21548
rect 10134 21536 10140 21548
rect 10095 21508 10140 21536
rect 10134 21496 10140 21508
rect 10192 21496 10198 21548
rect 12158 21536 12164 21548
rect 12119 21508 12164 21536
rect 12158 21496 12164 21508
rect 12216 21496 12222 21548
rect 14366 21496 14372 21548
rect 14424 21536 14430 21548
rect 14645 21539 14703 21545
rect 14645 21536 14657 21539
rect 14424 21508 14657 21536
rect 14424 21496 14430 21508
rect 14645 21505 14657 21508
rect 14691 21505 14703 21539
rect 15838 21536 15844 21548
rect 15799 21508 15844 21536
rect 14645 21499 14703 21505
rect 15838 21496 15844 21508
rect 15896 21496 15902 21548
rect 17313 21539 17371 21545
rect 17313 21505 17325 21539
rect 17359 21536 17371 21539
rect 17512 21536 17540 21564
rect 17770 21536 17776 21548
rect 17359 21508 17776 21536
rect 17359 21505 17371 21508
rect 17313 21499 17371 21505
rect 17770 21496 17776 21508
rect 17828 21496 17834 21548
rect 19996 21545 20024 21576
rect 26970 21564 26976 21616
rect 27028 21604 27034 21616
rect 29365 21607 29423 21613
rect 27028 21576 27922 21604
rect 27028 21564 27034 21576
rect 29365 21573 29377 21607
rect 29411 21604 29423 21607
rect 29730 21604 29736 21616
rect 29411 21576 29736 21604
rect 29411 21573 29423 21576
rect 29365 21567 29423 21573
rect 29730 21564 29736 21576
rect 29788 21564 29794 21616
rect 30374 21604 30380 21616
rect 30024 21576 30380 21604
rect 19981 21539 20039 21545
rect 19981 21505 19993 21539
rect 20027 21505 20039 21539
rect 19981 21499 20039 21505
rect 20809 21539 20867 21545
rect 20809 21505 20821 21539
rect 20855 21536 20867 21539
rect 21082 21536 21088 21548
rect 20855 21508 21088 21536
rect 20855 21505 20867 21508
rect 20809 21499 20867 21505
rect 21082 21496 21088 21508
rect 21140 21496 21146 21548
rect 22373 21539 22431 21545
rect 22373 21505 22385 21539
rect 22419 21536 22431 21539
rect 23566 21536 23572 21548
rect 22419 21508 23428 21536
rect 23527 21508 23572 21536
rect 22419 21505 22431 21508
rect 22373 21499 22431 21505
rect 13262 21468 13268 21480
rect 13175 21440 13268 21468
rect 13262 21428 13268 21440
rect 13320 21428 13326 21480
rect 13446 21468 13452 21480
rect 13407 21440 13452 21468
rect 13446 21428 13452 21440
rect 13504 21428 13510 21480
rect 16117 21471 16175 21477
rect 16117 21437 16129 21471
rect 16163 21468 16175 21471
rect 16482 21468 16488 21480
rect 16163 21440 16488 21468
rect 16163 21437 16175 21440
rect 16117 21431 16175 21437
rect 16482 21428 16488 21440
rect 16540 21428 16546 21480
rect 17589 21471 17647 21477
rect 17589 21437 17601 21471
rect 17635 21468 17647 21471
rect 17954 21468 17960 21480
rect 17635 21440 17960 21468
rect 17635 21437 17647 21440
rect 17589 21431 17647 21437
rect 17954 21428 17960 21440
rect 18012 21468 18018 21480
rect 18230 21468 18236 21480
rect 18012 21440 18236 21468
rect 18012 21428 18018 21440
rect 18230 21428 18236 21440
rect 18288 21428 18294 21480
rect 19702 21468 19708 21480
rect 19663 21440 19708 21468
rect 19702 21428 19708 21440
rect 19760 21428 19766 21480
rect 20990 21428 20996 21480
rect 21048 21468 21054 21480
rect 21048 21440 21093 21468
rect 21048 21428 21054 21440
rect 21818 21428 21824 21480
rect 21876 21468 21882 21480
rect 22557 21471 22615 21477
rect 21876 21440 22324 21468
rect 21876 21428 21882 21440
rect 13280 21400 13308 21428
rect 14734 21400 14740 21412
rect 13280 21372 14740 21400
rect 14734 21360 14740 21372
rect 14792 21360 14798 21412
rect 21910 21360 21916 21412
rect 21968 21400 21974 21412
rect 22005 21403 22063 21409
rect 22005 21400 22017 21403
rect 21968 21372 22017 21400
rect 21968 21360 21974 21372
rect 22005 21369 22017 21372
rect 22051 21369 22063 21403
rect 22296 21400 22324 21440
rect 22557 21437 22569 21471
rect 22603 21437 22615 21471
rect 22557 21431 22615 21437
rect 22572 21400 22600 21431
rect 22296 21372 22600 21400
rect 23400 21400 23428 21508
rect 23566 21496 23572 21508
rect 23624 21536 23630 21548
rect 24397 21539 24455 21545
rect 24397 21536 24409 21539
rect 23624 21508 24409 21536
rect 23624 21496 23630 21508
rect 24397 21505 24409 21508
rect 24443 21536 24455 21539
rect 24486 21536 24492 21548
rect 24443 21508 24492 21536
rect 24443 21505 24455 21508
rect 24397 21499 24455 21505
rect 24486 21496 24492 21508
rect 24544 21496 24550 21548
rect 26421 21539 26479 21545
rect 26421 21505 26433 21539
rect 26467 21536 26479 21539
rect 26510 21536 26516 21548
rect 26467 21508 26516 21536
rect 26467 21505 26479 21508
rect 26421 21499 26479 21505
rect 26510 21496 26516 21508
rect 26568 21496 26574 21548
rect 27154 21536 27160 21548
rect 27115 21508 27160 21536
rect 27154 21496 27160 21508
rect 27212 21496 27218 21548
rect 29641 21539 29699 21545
rect 29641 21505 29653 21539
rect 29687 21536 29699 21539
rect 30024 21536 30052 21576
rect 30374 21564 30380 21576
rect 30432 21564 30438 21616
rect 33502 21604 33508 21616
rect 32508 21576 33508 21604
rect 32508 21548 32536 21576
rect 33502 21564 33508 21576
rect 33560 21564 33566 21616
rect 35986 21564 35992 21616
rect 36044 21564 36050 21616
rect 30558 21536 30564 21548
rect 29687 21508 30052 21536
rect 30392 21508 30564 21536
rect 29687 21505 29699 21508
rect 29641 21499 29699 21505
rect 25590 21428 25596 21480
rect 25648 21468 25654 21480
rect 25774 21468 25780 21480
rect 25648 21440 25780 21468
rect 25648 21428 25654 21440
rect 25774 21428 25780 21440
rect 25832 21428 25838 21480
rect 30392 21477 30420 21508
rect 30558 21496 30564 21508
rect 30616 21496 30622 21548
rect 32490 21536 32496 21548
rect 31726 21508 32496 21536
rect 27433 21471 27491 21477
rect 27433 21468 27445 21471
rect 26620 21440 27445 21468
rect 26620 21409 26648 21440
rect 27433 21437 27445 21440
rect 27479 21437 27491 21471
rect 27433 21431 27491 21437
rect 30285 21471 30343 21477
rect 30285 21437 30297 21471
rect 30331 21437 30343 21471
rect 30285 21431 30343 21437
rect 30377 21471 30435 21477
rect 30377 21437 30389 21471
rect 30423 21437 30435 21471
rect 30377 21431 30435 21437
rect 26605 21403 26663 21409
rect 23400 21372 26556 21400
rect 22005 21363 22063 21369
rect 7834 21292 7840 21344
rect 7892 21332 7898 21344
rect 7929 21335 7987 21341
rect 7929 21332 7941 21335
rect 7892 21304 7941 21332
rect 7892 21292 7898 21304
rect 7929 21301 7941 21304
rect 7975 21301 7987 21335
rect 9950 21332 9956 21344
rect 9911 21304 9956 21332
rect 7929 21295 7987 21301
rect 9950 21292 9956 21304
rect 10008 21292 10014 21344
rect 16482 21292 16488 21344
rect 16540 21332 16546 21344
rect 18690 21332 18696 21344
rect 16540 21304 18696 21332
rect 16540 21292 16546 21304
rect 18690 21292 18696 21304
rect 18748 21292 18754 21344
rect 24302 21332 24308 21344
rect 24263 21304 24308 21332
rect 24302 21292 24308 21304
rect 24360 21292 24366 21344
rect 24946 21292 24952 21344
rect 25004 21332 25010 21344
rect 25225 21335 25283 21341
rect 25225 21332 25237 21335
rect 25004 21304 25237 21332
rect 25004 21292 25010 21304
rect 25225 21301 25237 21304
rect 25271 21301 25283 21335
rect 26528 21332 26556 21372
rect 26605 21369 26617 21403
rect 26651 21369 26663 21403
rect 29362 21400 29368 21412
rect 29323 21372 29368 21400
rect 26605 21363 26663 21369
rect 29362 21360 29368 21372
rect 29420 21360 29426 21412
rect 30300 21400 30328 21431
rect 30466 21428 30472 21480
rect 30524 21468 30530 21480
rect 31726 21468 31754 21508
rect 32490 21496 32496 21508
rect 32548 21496 32554 21548
rect 32582 21496 32588 21548
rect 32640 21536 32646 21548
rect 33781 21539 33839 21545
rect 33781 21536 33793 21539
rect 32640 21508 33793 21536
rect 32640 21496 32646 21508
rect 33781 21505 33793 21508
rect 33827 21505 33839 21539
rect 33781 21499 33839 21505
rect 32398 21468 32404 21480
rect 30524 21440 31754 21468
rect 32359 21440 32404 21468
rect 30524 21428 30530 21440
rect 32398 21428 32404 21440
rect 32456 21428 32462 21480
rect 33686 21468 33692 21480
rect 33647 21440 33692 21468
rect 33686 21428 33692 21440
rect 33744 21428 33750 21480
rect 34330 21428 34336 21480
rect 34388 21468 34394 21480
rect 34977 21471 35035 21477
rect 34977 21468 34989 21471
rect 34388 21440 34989 21468
rect 34388 21428 34394 21440
rect 34977 21437 34989 21440
rect 35023 21437 35035 21471
rect 34977 21431 35035 21437
rect 35253 21471 35311 21477
rect 35253 21437 35265 21471
rect 35299 21468 35311 21471
rect 35342 21468 35348 21480
rect 35299 21440 35348 21468
rect 35299 21437 35311 21440
rect 35253 21431 35311 21437
rect 35342 21428 35348 21440
rect 35400 21428 35406 21480
rect 31478 21400 31484 21412
rect 30300 21372 31484 21400
rect 30392 21344 30420 21372
rect 31478 21360 31484 21372
rect 31536 21360 31542 21412
rect 28626 21332 28632 21344
rect 26528 21304 28632 21332
rect 25225 21295 25283 21301
rect 28626 21292 28632 21304
rect 28684 21332 28690 21344
rect 30282 21332 30288 21344
rect 28684 21304 30288 21332
rect 28684 21292 28690 21304
rect 30282 21292 30288 21304
rect 30340 21292 30346 21344
rect 30374 21292 30380 21344
rect 30432 21292 30438 21344
rect 30834 21332 30840 21344
rect 30795 21304 30840 21332
rect 30834 21292 30840 21304
rect 30892 21292 30898 21344
rect 34054 21332 34060 21344
rect 34015 21304 34060 21332
rect 34054 21292 34060 21304
rect 34112 21292 34118 21344
rect 34790 21292 34796 21344
rect 34848 21332 34854 21344
rect 36725 21335 36783 21341
rect 36725 21332 36737 21335
rect 34848 21304 36737 21332
rect 34848 21292 34854 21304
rect 36725 21301 36737 21304
rect 36771 21301 36783 21335
rect 36725 21295 36783 21301
rect 1104 21242 37628 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 37628 21242
rect 1104 21168 37628 21190
rect 8570 21128 8576 21140
rect 8531 21100 8576 21128
rect 8570 21088 8576 21100
rect 8628 21088 8634 21140
rect 15838 21088 15844 21140
rect 15896 21128 15902 21140
rect 26510 21128 26516 21140
rect 15896 21100 22094 21128
rect 26471 21100 26516 21128
rect 15896 21088 15902 21100
rect 9582 21020 9588 21072
rect 9640 21020 9646 21072
rect 11974 21020 11980 21072
rect 12032 21060 12038 21072
rect 12526 21060 12532 21072
rect 12032 21032 12532 21060
rect 12032 21020 12038 21032
rect 12526 21020 12532 21032
rect 12584 21060 12590 21072
rect 22066 21060 22094 21100
rect 26510 21088 26516 21100
rect 26568 21088 26574 21140
rect 28718 21128 28724 21140
rect 28679 21100 28724 21128
rect 28718 21088 28724 21100
rect 28776 21088 28782 21140
rect 32398 21128 32404 21140
rect 30116 21100 32404 21128
rect 26786 21060 26792 21072
rect 12584 21032 16436 21060
rect 22066 21032 26792 21060
rect 12584 21020 12590 21032
rect 6822 20992 6828 21004
rect 6783 20964 6828 20992
rect 6822 20952 6828 20964
rect 6880 20952 6886 21004
rect 9600 20992 9628 21020
rect 9677 20995 9735 21001
rect 9677 20992 9689 20995
rect 9600 20964 9689 20992
rect 9677 20961 9689 20964
rect 9723 20961 9735 20995
rect 9677 20955 9735 20961
rect 10870 20952 10876 21004
rect 10928 20992 10934 21004
rect 12618 20992 12624 21004
rect 10928 20964 12296 20992
rect 12579 20964 12624 20992
rect 10928 20952 10934 20964
rect 9493 20927 9551 20933
rect 9493 20893 9505 20927
rect 9539 20924 9551 20927
rect 9582 20924 9588 20936
rect 9539 20896 9588 20924
rect 9539 20893 9551 20896
rect 9493 20887 9551 20893
rect 9582 20884 9588 20896
rect 9640 20884 9646 20936
rect 10980 20933 11008 20964
rect 10965 20927 11023 20933
rect 10965 20893 10977 20927
rect 11011 20893 11023 20927
rect 10965 20887 11023 20893
rect 11425 20927 11483 20933
rect 11425 20893 11437 20927
rect 11471 20924 11483 20927
rect 11471 20896 12112 20924
rect 11471 20893 11483 20896
rect 11425 20887 11483 20893
rect 7098 20856 7104 20868
rect 7059 20828 7104 20856
rect 7098 20816 7104 20828
rect 7156 20816 7162 20868
rect 7834 20816 7840 20868
rect 7892 20816 7898 20868
rect 8754 20816 8760 20868
rect 8812 20856 8818 20868
rect 8812 20828 9628 20856
rect 8812 20816 8818 20828
rect 8662 20748 8668 20800
rect 8720 20788 8726 20800
rect 9600 20797 9628 20828
rect 9125 20791 9183 20797
rect 9125 20788 9137 20791
rect 8720 20760 9137 20788
rect 8720 20748 8726 20760
rect 9125 20757 9137 20760
rect 9171 20757 9183 20791
rect 9125 20751 9183 20757
rect 9585 20791 9643 20797
rect 9585 20757 9597 20791
rect 9631 20757 9643 20791
rect 9585 20751 9643 20757
rect 10778 20748 10784 20800
rect 10836 20788 10842 20800
rect 10873 20791 10931 20797
rect 10873 20788 10885 20791
rect 10836 20760 10885 20788
rect 10836 20748 10842 20760
rect 10873 20757 10885 20760
rect 10919 20757 10931 20791
rect 11606 20788 11612 20800
rect 11567 20760 11612 20788
rect 10873 20751 10931 20757
rect 11606 20748 11612 20760
rect 11664 20748 11670 20800
rect 12084 20797 12112 20896
rect 12268 20856 12296 20964
rect 12618 20952 12624 20964
rect 12676 20952 12682 21004
rect 16408 20992 16436 21032
rect 26786 21020 26792 21032
rect 26844 21060 26850 21072
rect 26844 21032 27292 21060
rect 26844 21020 26850 21032
rect 19613 20995 19671 21001
rect 19613 20992 19625 20995
rect 16408 20964 19625 20992
rect 19613 20961 19625 20964
rect 19659 20992 19671 20995
rect 20070 20992 20076 21004
rect 19659 20964 20076 20992
rect 19659 20961 19671 20964
rect 19613 20955 19671 20961
rect 20070 20952 20076 20964
rect 20128 20952 20134 21004
rect 20714 20952 20720 21004
rect 20772 20992 20778 21004
rect 21818 20992 21824 21004
rect 20772 20964 21824 20992
rect 20772 20952 20778 20964
rect 21818 20952 21824 20964
rect 21876 20992 21882 21004
rect 22373 20995 22431 21001
rect 22373 20992 22385 20995
rect 21876 20964 22385 20992
rect 21876 20952 21882 20964
rect 22373 20961 22385 20964
rect 22419 20961 22431 20995
rect 22373 20955 22431 20961
rect 23293 20995 23351 21001
rect 23293 20961 23305 20995
rect 23339 20992 23351 20995
rect 23566 20992 23572 21004
rect 23339 20964 23572 20992
rect 23339 20961 23351 20964
rect 23293 20955 23351 20961
rect 23566 20952 23572 20964
rect 23624 20952 23630 21004
rect 25130 20992 25136 21004
rect 25091 20964 25136 20992
rect 25130 20952 25136 20964
rect 25188 20952 25194 21004
rect 25314 20952 25320 21004
rect 25372 20992 25378 21004
rect 25682 20992 25688 21004
rect 25372 20964 25688 20992
rect 25372 20952 25378 20964
rect 25682 20952 25688 20964
rect 25740 20992 25746 21004
rect 25869 20995 25927 21001
rect 25869 20992 25881 20995
rect 25740 20964 25881 20992
rect 25740 20952 25746 20964
rect 25869 20961 25881 20964
rect 25915 20961 25927 20995
rect 25869 20955 25927 20961
rect 27264 20992 27292 21032
rect 27522 20992 27528 21004
rect 27264 20964 27528 20992
rect 12434 20884 12440 20936
rect 12492 20924 12498 20936
rect 14274 20924 14280 20936
rect 12492 20896 12537 20924
rect 14235 20896 14280 20924
rect 12492 20884 12498 20896
rect 14274 20884 14280 20896
rect 14332 20884 14338 20936
rect 14366 20884 14372 20936
rect 14424 20924 14430 20936
rect 15381 20927 15439 20933
rect 15381 20924 15393 20927
rect 14424 20896 15393 20924
rect 14424 20884 14430 20896
rect 15381 20893 15393 20896
rect 15427 20893 15439 20927
rect 15381 20887 15439 20893
rect 17678 20884 17684 20936
rect 17736 20924 17742 20936
rect 19886 20924 19892 20936
rect 17736 20896 19892 20924
rect 17736 20884 17742 20896
rect 19886 20884 19892 20896
rect 19944 20884 19950 20936
rect 23017 20927 23075 20933
rect 23017 20924 23029 20927
rect 22112 20896 23029 20924
rect 14384 20856 14412 20884
rect 22112 20868 22140 20896
rect 23017 20893 23029 20896
rect 23063 20893 23075 20927
rect 24946 20924 24952 20936
rect 24907 20896 24952 20924
rect 23017 20887 23075 20893
rect 24946 20884 24952 20896
rect 25004 20884 25010 20936
rect 27264 20933 27292 20964
rect 27522 20952 27528 20964
rect 27580 20952 27586 21004
rect 29089 20995 29147 21001
rect 29089 20961 29101 20995
rect 29135 20992 29147 20995
rect 30116 20992 30144 21100
rect 32398 21088 32404 21100
rect 32456 21088 32462 21140
rect 32953 21131 33011 21137
rect 32953 21097 32965 21131
rect 32999 21128 33011 21131
rect 33686 21128 33692 21140
rect 32999 21100 33692 21128
rect 32999 21097 33011 21100
rect 32953 21091 33011 21097
rect 33686 21088 33692 21100
rect 33744 21088 33750 21140
rect 31478 21020 31484 21072
rect 31536 21060 31542 21072
rect 34606 21060 34612 21072
rect 31536 21032 34612 21060
rect 31536 21020 31542 21032
rect 29135 20964 30144 20992
rect 30193 20995 30251 21001
rect 29135 20961 29147 20964
rect 29089 20955 29147 20961
rect 30193 20961 30205 20995
rect 30239 20992 30251 20995
rect 31202 20992 31208 21004
rect 30239 20964 31208 20992
rect 30239 20961 30251 20964
rect 30193 20955 30251 20961
rect 31202 20952 31208 20964
rect 31260 20952 31266 21004
rect 33520 21001 33548 21032
rect 34606 21020 34612 21032
rect 34664 21060 34670 21072
rect 34664 21032 35480 21060
rect 34664 21020 34670 21032
rect 33505 20995 33563 21001
rect 33505 20961 33517 20995
rect 33551 20961 33563 20995
rect 33505 20955 33563 20961
rect 34790 20952 34796 21004
rect 34848 20992 34854 21004
rect 35452 21001 35480 21032
rect 35345 20995 35403 21001
rect 35345 20992 35357 20995
rect 34848 20964 35357 20992
rect 34848 20952 34854 20964
rect 35345 20961 35357 20964
rect 35391 20961 35403 20995
rect 35345 20955 35403 20961
rect 35437 20995 35495 21001
rect 35437 20961 35449 20995
rect 35483 20961 35495 20995
rect 35437 20955 35495 20961
rect 27249 20927 27307 20933
rect 27249 20893 27261 20927
rect 27295 20893 27307 20927
rect 28442 20924 28448 20936
rect 27249 20887 27307 20893
rect 27356 20896 28448 20924
rect 12268 20828 14412 20856
rect 16666 20816 16672 20868
rect 16724 20816 16730 20868
rect 17402 20856 17408 20868
rect 17363 20828 17408 20856
rect 17402 20816 17408 20828
rect 17460 20816 17466 20868
rect 18046 20816 18052 20868
rect 18104 20856 18110 20868
rect 18506 20856 18512 20868
rect 18104 20828 18512 20856
rect 18104 20816 18110 20828
rect 18506 20816 18512 20828
rect 18564 20816 18570 20868
rect 21358 20856 21364 20868
rect 21319 20828 21364 20856
rect 21358 20816 21364 20828
rect 21416 20816 21422 20868
rect 22094 20856 22100 20868
rect 21468 20828 22100 20856
rect 12069 20791 12127 20797
rect 12069 20757 12081 20791
rect 12115 20757 12127 20791
rect 12069 20751 12127 20757
rect 12529 20791 12587 20797
rect 12529 20757 12541 20791
rect 12575 20788 12587 20791
rect 13446 20788 13452 20800
rect 12575 20760 13452 20788
rect 12575 20757 12587 20760
rect 12529 20751 12587 20757
rect 13446 20748 13452 20760
rect 13504 20748 13510 20800
rect 14458 20788 14464 20800
rect 14419 20760 14464 20788
rect 14458 20748 14464 20760
rect 14516 20748 14522 20800
rect 15289 20791 15347 20797
rect 15289 20757 15301 20791
rect 15335 20788 15347 20791
rect 15378 20788 15384 20800
rect 15335 20760 15384 20788
rect 15335 20757 15347 20760
rect 15289 20751 15347 20757
rect 15378 20748 15384 20760
rect 15436 20748 15442 20800
rect 15654 20748 15660 20800
rect 15712 20788 15718 20800
rect 15933 20791 15991 20797
rect 15933 20788 15945 20791
rect 15712 20760 15945 20788
rect 15712 20748 15718 20760
rect 15933 20757 15945 20760
rect 15979 20757 15991 20791
rect 15933 20751 15991 20757
rect 17770 20748 17776 20800
rect 17828 20788 17834 20800
rect 18785 20791 18843 20797
rect 18785 20788 18797 20791
rect 17828 20760 18797 20788
rect 17828 20748 17834 20760
rect 18785 20757 18797 20760
rect 18831 20788 18843 20791
rect 21468 20788 21496 20828
rect 22094 20816 22100 20828
rect 22152 20816 22158 20868
rect 22189 20859 22247 20865
rect 22189 20825 22201 20859
rect 22235 20856 22247 20859
rect 27356 20856 27384 20896
rect 28442 20884 28448 20896
rect 28500 20884 28506 20936
rect 28994 20924 29000 20936
rect 28907 20896 29000 20924
rect 28994 20884 29000 20896
rect 29052 20924 29058 20936
rect 29730 20924 29736 20936
rect 29052 20896 29736 20924
rect 29052 20884 29058 20896
rect 29730 20884 29736 20896
rect 29788 20884 29794 20936
rect 31570 20884 31576 20936
rect 31628 20884 31634 20936
rect 32677 20927 32735 20933
rect 32677 20893 32689 20927
rect 32723 20893 32735 20927
rect 32677 20887 32735 20893
rect 32769 20927 32827 20933
rect 32769 20893 32781 20927
rect 32815 20924 32827 20927
rect 32858 20924 32864 20936
rect 32815 20896 32864 20924
rect 32815 20893 32827 20896
rect 32769 20887 32827 20893
rect 22235 20828 27384 20856
rect 27525 20859 27583 20865
rect 22235 20825 22247 20828
rect 22189 20819 22247 20825
rect 27525 20825 27537 20859
rect 27571 20856 27583 20859
rect 27706 20856 27712 20868
rect 27571 20828 27712 20856
rect 27571 20825 27583 20828
rect 27525 20819 27583 20825
rect 27706 20816 27712 20828
rect 27764 20856 27770 20868
rect 28718 20856 28724 20868
rect 27764 20828 28724 20856
rect 27764 20816 27770 20828
rect 28718 20816 28724 20828
rect 28776 20816 28782 20868
rect 30466 20856 30472 20868
rect 30427 20828 30472 20856
rect 30466 20816 30472 20828
rect 30524 20816 30530 20868
rect 32692 20856 32720 20887
rect 32858 20884 32864 20896
rect 32916 20884 32922 20936
rect 32953 20927 33011 20933
rect 32953 20893 32965 20927
rect 32999 20924 33011 20927
rect 33594 20924 33600 20936
rect 32999 20896 33600 20924
rect 32999 20893 33011 20896
rect 32953 20887 33011 20893
rect 33594 20884 33600 20896
rect 33652 20884 33658 20936
rect 34054 20884 34060 20936
rect 34112 20924 34118 20936
rect 35253 20927 35311 20933
rect 35253 20924 35265 20927
rect 34112 20896 35265 20924
rect 34112 20884 34118 20896
rect 35253 20893 35265 20896
rect 35299 20893 35311 20927
rect 35253 20887 35311 20893
rect 33410 20856 33416 20868
rect 32692 20828 33416 20856
rect 33410 20816 33416 20828
rect 33468 20816 33474 20868
rect 33502 20816 33508 20868
rect 33560 20856 33566 20868
rect 33689 20859 33747 20865
rect 33689 20856 33701 20859
rect 33560 20828 33701 20856
rect 33560 20816 33566 20828
rect 33689 20825 33701 20828
rect 33735 20825 33747 20859
rect 33689 20819 33747 20825
rect 21818 20788 21824 20800
rect 18831 20760 21496 20788
rect 21779 20760 21824 20788
rect 18831 20757 18843 20760
rect 18785 20751 18843 20757
rect 21818 20748 21824 20760
rect 21876 20748 21882 20800
rect 22278 20748 22284 20800
rect 22336 20788 22342 20800
rect 24581 20791 24639 20797
rect 22336 20760 22381 20788
rect 22336 20748 22342 20760
rect 24581 20757 24593 20791
rect 24627 20788 24639 20791
rect 24762 20788 24768 20800
rect 24627 20760 24768 20788
rect 24627 20757 24639 20760
rect 24581 20751 24639 20757
rect 24762 20748 24768 20760
rect 24820 20748 24826 20800
rect 25041 20791 25099 20797
rect 25041 20757 25053 20791
rect 25087 20788 25099 20791
rect 25590 20788 25596 20800
rect 25087 20760 25596 20788
rect 25087 20757 25099 20760
rect 25041 20751 25099 20757
rect 25590 20748 25596 20760
rect 25648 20788 25654 20800
rect 26053 20791 26111 20797
rect 26053 20788 26065 20791
rect 25648 20760 26065 20788
rect 25648 20748 25654 20760
rect 26053 20757 26065 20760
rect 26099 20757 26111 20791
rect 26053 20751 26111 20757
rect 26145 20791 26203 20797
rect 26145 20757 26157 20791
rect 26191 20788 26203 20791
rect 27246 20788 27252 20800
rect 26191 20760 27252 20788
rect 26191 20757 26203 20760
rect 26145 20751 26203 20757
rect 27246 20748 27252 20760
rect 27304 20748 27310 20800
rect 30558 20748 30564 20800
rect 30616 20788 30622 20800
rect 31941 20791 31999 20797
rect 31941 20788 31953 20791
rect 30616 20760 31953 20788
rect 30616 20748 30622 20760
rect 31941 20757 31953 20760
rect 31987 20757 31999 20791
rect 31941 20751 31999 20757
rect 33778 20748 33784 20800
rect 33836 20788 33842 20800
rect 34146 20788 34152 20800
rect 33836 20760 33881 20788
rect 34107 20760 34152 20788
rect 33836 20748 33842 20760
rect 34146 20748 34152 20760
rect 34204 20748 34210 20800
rect 34885 20791 34943 20797
rect 34885 20757 34897 20791
rect 34931 20788 34943 20791
rect 34974 20788 34980 20800
rect 34931 20760 34980 20788
rect 34931 20757 34943 20760
rect 34885 20751 34943 20757
rect 34974 20748 34980 20760
rect 35032 20748 35038 20800
rect 1104 20698 37628 20720
rect 1104 20646 4874 20698
rect 4926 20646 4938 20698
rect 4990 20646 5002 20698
rect 5054 20646 5066 20698
rect 5118 20646 5130 20698
rect 5182 20646 35594 20698
rect 35646 20646 35658 20698
rect 35710 20646 35722 20698
rect 35774 20646 35786 20698
rect 35838 20646 35850 20698
rect 35902 20646 37628 20698
rect 1104 20624 37628 20646
rect 7098 20544 7104 20596
rect 7156 20584 7162 20596
rect 7377 20587 7435 20593
rect 7377 20584 7389 20587
rect 7156 20556 7389 20584
rect 7156 20544 7162 20556
rect 7377 20553 7389 20556
rect 7423 20553 7435 20587
rect 7377 20547 7435 20553
rect 8389 20587 8447 20593
rect 8389 20553 8401 20587
rect 8435 20584 8447 20587
rect 8662 20584 8668 20596
rect 8435 20556 8668 20584
rect 8435 20553 8447 20556
rect 8389 20547 8447 20553
rect 8662 20544 8668 20556
rect 8720 20544 8726 20596
rect 11149 20587 11207 20593
rect 11149 20553 11161 20587
rect 11195 20584 11207 20587
rect 11514 20584 11520 20596
rect 11195 20556 11520 20584
rect 11195 20553 11207 20556
rect 11149 20547 11207 20553
rect 11514 20544 11520 20556
rect 11572 20584 11578 20596
rect 12894 20584 12900 20596
rect 11572 20556 12900 20584
rect 11572 20544 11578 20556
rect 12894 20544 12900 20556
rect 12952 20584 12958 20596
rect 13446 20584 13452 20596
rect 12952 20556 13308 20584
rect 13407 20556 13452 20584
rect 12952 20544 12958 20556
rect 6822 20476 6828 20528
rect 6880 20516 6886 20528
rect 8294 20516 8300 20528
rect 6880 20488 8300 20516
rect 6880 20476 6886 20488
rect 8294 20476 8300 20488
rect 8352 20516 8358 20528
rect 9677 20519 9735 20525
rect 8352 20488 9168 20516
rect 8352 20476 8358 20488
rect 9140 20460 9168 20488
rect 9677 20485 9689 20519
rect 9723 20516 9735 20519
rect 9950 20516 9956 20528
rect 9723 20488 9956 20516
rect 9723 20485 9735 20488
rect 9677 20479 9735 20485
rect 9950 20476 9956 20488
rect 10008 20476 10014 20528
rect 11606 20476 11612 20528
rect 11664 20516 11670 20528
rect 11977 20519 12035 20525
rect 11977 20516 11989 20519
rect 11664 20488 11989 20516
rect 11664 20476 11670 20488
rect 11977 20485 11989 20488
rect 12023 20485 12035 20519
rect 11977 20479 12035 20485
rect 12434 20476 12440 20528
rect 12492 20476 12498 20528
rect 13280 20516 13308 20556
rect 13446 20544 13452 20556
rect 13504 20544 13510 20596
rect 15654 20584 15660 20596
rect 13556 20556 15660 20584
rect 13556 20516 13584 20556
rect 15654 20544 15660 20556
rect 15712 20544 15718 20596
rect 15841 20587 15899 20593
rect 15841 20553 15853 20587
rect 15887 20584 15899 20587
rect 15930 20584 15936 20596
rect 15887 20556 15936 20584
rect 15887 20553 15899 20556
rect 15841 20547 15899 20553
rect 15930 20544 15936 20556
rect 15988 20544 15994 20596
rect 17037 20587 17095 20593
rect 17037 20553 17049 20587
rect 17083 20584 17095 20587
rect 17402 20584 17408 20596
rect 17083 20556 17408 20584
rect 17083 20553 17095 20556
rect 17037 20547 17095 20553
rect 17402 20544 17408 20556
rect 17460 20544 17466 20596
rect 19426 20544 19432 20596
rect 19484 20584 19490 20596
rect 19705 20587 19763 20593
rect 19705 20584 19717 20587
rect 19484 20556 19717 20584
rect 19484 20544 19490 20556
rect 19705 20553 19717 20556
rect 19751 20553 19763 20587
rect 19705 20547 19763 20553
rect 24765 20587 24823 20593
rect 24765 20553 24777 20587
rect 24811 20584 24823 20587
rect 25590 20584 25596 20596
rect 24811 20556 25596 20584
rect 24811 20553 24823 20556
rect 24765 20547 24823 20553
rect 25590 20544 25596 20556
rect 25648 20544 25654 20596
rect 25685 20587 25743 20593
rect 25685 20553 25697 20587
rect 25731 20584 25743 20587
rect 27525 20587 27583 20593
rect 27525 20584 27537 20587
rect 25731 20556 27537 20584
rect 25731 20553 25743 20556
rect 25685 20547 25743 20553
rect 27525 20553 27537 20556
rect 27571 20584 27583 20587
rect 28166 20584 28172 20596
rect 27571 20556 28172 20584
rect 27571 20553 27583 20556
rect 27525 20547 27583 20553
rect 28166 20544 28172 20556
rect 28224 20544 28230 20596
rect 29178 20544 29184 20596
rect 29236 20584 29242 20596
rect 29825 20587 29883 20593
rect 29825 20584 29837 20587
rect 29236 20556 29837 20584
rect 29236 20544 29242 20556
rect 29825 20553 29837 20556
rect 29871 20553 29883 20587
rect 29825 20547 29883 20553
rect 30193 20587 30251 20593
rect 30193 20553 30205 20587
rect 30239 20553 30251 20587
rect 30193 20547 30251 20553
rect 13280 20488 13584 20516
rect 14369 20519 14427 20525
rect 14369 20485 14381 20519
rect 14415 20516 14427 20519
rect 14458 20516 14464 20528
rect 14415 20488 14464 20516
rect 14415 20485 14427 20488
rect 14369 20479 14427 20485
rect 14458 20476 14464 20488
rect 14516 20476 14522 20528
rect 15378 20476 15384 20528
rect 15436 20476 15442 20528
rect 21818 20516 21824 20528
rect 16868 20488 21824 20516
rect 1765 20451 1823 20457
rect 1765 20417 1777 20451
rect 1811 20448 1823 20451
rect 2130 20448 2136 20460
rect 1811 20420 2136 20448
rect 1811 20417 1823 20420
rect 1765 20411 1823 20417
rect 2130 20408 2136 20420
rect 2188 20408 2194 20460
rect 7561 20451 7619 20457
rect 7561 20417 7573 20451
rect 7607 20448 7619 20451
rect 8478 20448 8484 20460
rect 7607 20420 8064 20448
rect 8439 20420 8484 20448
rect 7607 20417 7619 20420
rect 7561 20411 7619 20417
rect 1578 20312 1584 20324
rect 1539 20284 1584 20312
rect 1578 20272 1584 20284
rect 1636 20272 1642 20324
rect 8036 20321 8064 20420
rect 8478 20408 8484 20420
rect 8536 20408 8542 20460
rect 9122 20408 9128 20460
rect 9180 20448 9186 20460
rect 9401 20451 9459 20457
rect 9401 20448 9413 20451
rect 9180 20420 9413 20448
rect 9180 20408 9186 20420
rect 9401 20417 9413 20420
rect 9447 20417 9459 20451
rect 9401 20411 9459 20417
rect 10778 20408 10784 20460
rect 10836 20408 10842 20460
rect 11698 20448 11704 20460
rect 11659 20420 11704 20448
rect 11698 20408 11704 20420
rect 11756 20408 11762 20460
rect 16868 20457 16896 20488
rect 21818 20476 21824 20488
rect 21876 20476 21882 20528
rect 24670 20516 24676 20528
rect 24518 20488 24676 20516
rect 24670 20476 24676 20488
rect 24728 20476 24734 20528
rect 25314 20476 25320 20528
rect 25372 20516 25378 20528
rect 30208 20516 30236 20547
rect 30466 20544 30472 20596
rect 30524 20584 30530 20596
rect 30653 20587 30711 20593
rect 30653 20584 30665 20587
rect 30524 20556 30665 20584
rect 30524 20544 30530 20556
rect 30653 20553 30665 20556
rect 30699 20553 30711 20587
rect 30653 20547 30711 20553
rect 31570 20544 31576 20596
rect 31628 20584 31634 20596
rect 32401 20587 32459 20593
rect 32401 20584 32413 20587
rect 31628 20556 32413 20584
rect 31628 20544 31634 20556
rect 32401 20553 32413 20556
rect 32447 20553 32459 20587
rect 32401 20547 32459 20553
rect 35161 20587 35219 20593
rect 35161 20553 35173 20587
rect 35207 20584 35219 20587
rect 35342 20584 35348 20596
rect 35207 20556 35348 20584
rect 35207 20553 35219 20556
rect 35161 20547 35219 20553
rect 35342 20544 35348 20556
rect 35400 20544 35406 20596
rect 36078 20516 36084 20528
rect 25372 20488 27568 20516
rect 30208 20488 31524 20516
rect 25372 20476 25378 20488
rect 16853 20451 16911 20457
rect 16853 20417 16865 20451
rect 16899 20417 16911 20451
rect 16853 20411 16911 20417
rect 17681 20451 17739 20457
rect 17681 20417 17693 20451
rect 17727 20448 17739 20451
rect 17770 20448 17776 20460
rect 17727 20420 17776 20448
rect 17727 20417 17739 20420
rect 17681 20411 17739 20417
rect 17770 20408 17776 20420
rect 17828 20408 17834 20460
rect 18601 20451 18659 20457
rect 18601 20417 18613 20451
rect 18647 20448 18659 20451
rect 19613 20451 19671 20457
rect 18647 20420 19288 20448
rect 18647 20417 18659 20420
rect 18601 20411 18659 20417
rect 8665 20383 8723 20389
rect 8665 20349 8677 20383
rect 8711 20380 8723 20383
rect 10686 20380 10692 20392
rect 8711 20352 10692 20380
rect 8711 20349 8723 20352
rect 8665 20343 8723 20349
rect 10686 20340 10692 20352
rect 10744 20340 10750 20392
rect 14090 20380 14096 20392
rect 14051 20352 14096 20380
rect 14090 20340 14096 20352
rect 14148 20340 14154 20392
rect 19260 20321 19288 20420
rect 19613 20417 19625 20451
rect 19659 20417 19671 20451
rect 20622 20448 20628 20460
rect 20583 20420 20628 20448
rect 19613 20411 19671 20417
rect 8021 20315 8079 20321
rect 8021 20281 8033 20315
rect 8067 20281 8079 20315
rect 8021 20275 8079 20281
rect 19245 20315 19303 20321
rect 19245 20281 19257 20315
rect 19291 20281 19303 20315
rect 19628 20312 19656 20411
rect 20622 20408 20628 20420
rect 20680 20408 20686 20460
rect 21174 20408 21180 20460
rect 21232 20448 21238 20460
rect 21269 20451 21327 20457
rect 21269 20448 21281 20451
rect 21232 20420 21281 20448
rect 21232 20408 21238 20420
rect 21269 20417 21281 20420
rect 21315 20417 21327 20451
rect 22554 20448 22560 20460
rect 22515 20420 22560 20448
rect 21269 20411 21327 20417
rect 22554 20408 22560 20420
rect 22612 20408 22618 20460
rect 26421 20451 26479 20457
rect 26421 20417 26433 20451
rect 26467 20448 26479 20451
rect 27540 20448 27568 20488
rect 28537 20451 28595 20457
rect 26467 20420 27200 20448
rect 27540 20420 27752 20448
rect 26467 20417 26479 20420
rect 26421 20411 26479 20417
rect 19794 20380 19800 20392
rect 19755 20352 19800 20380
rect 19794 20340 19800 20352
rect 19852 20380 19858 20392
rect 20714 20380 20720 20392
rect 19852 20352 20720 20380
rect 19852 20340 19858 20352
rect 20714 20340 20720 20352
rect 20772 20340 20778 20392
rect 22002 20340 22008 20392
rect 22060 20380 22066 20392
rect 23017 20383 23075 20389
rect 23017 20380 23029 20383
rect 22060 20352 23029 20380
rect 22060 20340 22066 20352
rect 23017 20349 23029 20352
rect 23063 20349 23075 20383
rect 23017 20343 23075 20349
rect 23293 20383 23351 20389
rect 23293 20349 23305 20383
rect 23339 20380 23351 20383
rect 24578 20380 24584 20392
rect 23339 20352 24584 20380
rect 23339 20349 23351 20352
rect 23293 20343 23351 20349
rect 24578 20340 24584 20352
rect 24636 20340 24642 20392
rect 25774 20380 25780 20392
rect 25735 20352 25780 20380
rect 25774 20340 25780 20352
rect 25832 20340 25838 20392
rect 27172 20321 27200 20420
rect 27246 20340 27252 20392
rect 27304 20380 27310 20392
rect 27724 20389 27752 20420
rect 28537 20417 28549 20451
rect 28583 20448 28595 20451
rect 28718 20448 28724 20460
rect 28583 20420 28724 20448
rect 28583 20417 28595 20420
rect 28537 20411 28595 20417
rect 28718 20408 28724 20420
rect 28776 20408 28782 20460
rect 30374 20448 30380 20460
rect 29656 20420 30380 20448
rect 29656 20389 29684 20420
rect 30374 20408 30380 20420
rect 30432 20408 30438 20460
rect 30834 20448 30840 20460
rect 30795 20420 30840 20448
rect 30834 20408 30840 20420
rect 30892 20408 30898 20460
rect 31496 20457 31524 20488
rect 32508 20488 36084 20516
rect 31481 20451 31539 20457
rect 31481 20417 31493 20451
rect 31527 20417 31539 20451
rect 31481 20411 31539 20417
rect 31570 20408 31576 20460
rect 31628 20448 31634 20460
rect 32508 20457 32536 20488
rect 32493 20451 32551 20457
rect 32493 20448 32505 20451
rect 31628 20420 32505 20448
rect 31628 20408 31634 20420
rect 32493 20417 32505 20420
rect 32539 20417 32551 20451
rect 32493 20411 32551 20417
rect 32858 20408 32864 20460
rect 32916 20448 32922 20460
rect 33505 20451 33563 20457
rect 33505 20448 33517 20451
rect 32916 20420 33517 20448
rect 32916 20408 32922 20420
rect 33505 20417 33517 20420
rect 33551 20417 33563 20451
rect 33505 20411 33563 20417
rect 34146 20408 34152 20460
rect 34204 20448 34210 20460
rect 34517 20451 34575 20457
rect 34517 20448 34529 20451
rect 34204 20420 34529 20448
rect 34204 20408 34210 20420
rect 34517 20417 34529 20420
rect 34563 20417 34575 20451
rect 34974 20448 34980 20460
rect 34935 20420 34980 20448
rect 34517 20411 34575 20417
rect 34974 20408 34980 20420
rect 35032 20408 35038 20460
rect 35820 20457 35848 20488
rect 36078 20476 36084 20488
rect 36136 20476 36142 20528
rect 35805 20451 35863 20457
rect 35805 20417 35817 20451
rect 35851 20417 35863 20451
rect 35805 20411 35863 20417
rect 36630 20408 36636 20460
rect 36688 20448 36694 20460
rect 36725 20451 36783 20457
rect 36725 20448 36737 20451
rect 36688 20420 36737 20448
rect 36688 20408 36694 20420
rect 36725 20417 36737 20420
rect 36771 20417 36783 20451
rect 36725 20411 36783 20417
rect 27617 20383 27675 20389
rect 27617 20380 27629 20383
rect 27304 20352 27629 20380
rect 27304 20340 27310 20352
rect 27617 20349 27629 20352
rect 27663 20349 27675 20383
rect 27617 20343 27675 20349
rect 27709 20383 27767 20389
rect 27709 20349 27721 20383
rect 27755 20349 27767 20383
rect 27709 20343 27767 20349
rect 29641 20383 29699 20389
rect 29641 20349 29653 20383
rect 29687 20349 29699 20383
rect 29641 20343 29699 20349
rect 29730 20340 29736 20392
rect 29788 20380 29794 20392
rect 33410 20380 33416 20392
rect 29788 20352 29833 20380
rect 33371 20352 33416 20380
rect 29788 20340 29794 20352
rect 33410 20340 33416 20352
rect 33468 20340 33474 20392
rect 33778 20340 33784 20392
rect 33836 20380 33842 20392
rect 33873 20383 33931 20389
rect 33873 20380 33885 20383
rect 33836 20352 33885 20380
rect 33836 20340 33842 20352
rect 33873 20349 33885 20352
rect 33919 20349 33931 20383
rect 33873 20343 33931 20349
rect 27157 20315 27215 20321
rect 19628 20284 23152 20312
rect 19245 20275 19303 20281
rect 17586 20244 17592 20256
rect 17547 20216 17592 20244
rect 17586 20204 17592 20216
rect 17644 20204 17650 20256
rect 18785 20247 18843 20253
rect 18785 20213 18797 20247
rect 18831 20244 18843 20247
rect 19150 20244 19156 20256
rect 18831 20216 19156 20244
rect 18831 20213 18843 20216
rect 18785 20207 18843 20213
rect 19150 20204 19156 20216
rect 19208 20204 19214 20256
rect 20714 20204 20720 20256
rect 20772 20244 20778 20256
rect 20809 20247 20867 20253
rect 20809 20244 20821 20247
rect 20772 20216 20821 20244
rect 20772 20204 20778 20216
rect 20809 20213 20821 20216
rect 20855 20213 20867 20247
rect 20809 20207 20867 20213
rect 21266 20204 21272 20256
rect 21324 20244 21330 20256
rect 21361 20247 21419 20253
rect 21361 20244 21373 20247
rect 21324 20216 21373 20244
rect 21324 20204 21330 20216
rect 21361 20213 21373 20216
rect 21407 20213 21419 20247
rect 22370 20244 22376 20256
rect 22331 20216 22376 20244
rect 21361 20207 21419 20213
rect 22370 20204 22376 20216
rect 22428 20204 22434 20256
rect 23124 20244 23152 20284
rect 25056 20284 27108 20312
rect 25056 20244 25084 20284
rect 25222 20244 25228 20256
rect 23124 20216 25084 20244
rect 25183 20216 25228 20244
rect 25222 20204 25228 20216
rect 25280 20204 25286 20256
rect 26605 20247 26663 20253
rect 26605 20213 26617 20247
rect 26651 20244 26663 20247
rect 26970 20244 26976 20256
rect 26651 20216 26976 20244
rect 26651 20213 26663 20216
rect 26605 20207 26663 20213
rect 26970 20204 26976 20216
rect 27028 20204 27034 20256
rect 27080 20244 27108 20284
rect 27157 20281 27169 20315
rect 27203 20281 27215 20315
rect 30558 20312 30564 20324
rect 27157 20275 27215 20281
rect 28184 20284 30564 20312
rect 28184 20244 28212 20284
rect 30558 20272 30564 20284
rect 30616 20272 30622 20324
rect 36906 20312 36912 20324
rect 36867 20284 36912 20312
rect 36906 20272 36912 20284
rect 36964 20272 36970 20324
rect 27080 20216 28212 20244
rect 28258 20204 28264 20256
rect 28316 20244 28322 20256
rect 28445 20247 28503 20253
rect 28445 20244 28457 20247
rect 28316 20216 28457 20244
rect 28316 20204 28322 20216
rect 28445 20213 28457 20216
rect 28491 20213 28503 20247
rect 31294 20244 31300 20256
rect 31255 20216 31300 20244
rect 28445 20207 28503 20213
rect 31294 20204 31300 20216
rect 31352 20204 31358 20256
rect 34054 20204 34060 20256
rect 34112 20244 34118 20256
rect 34333 20247 34391 20253
rect 34333 20244 34345 20247
rect 34112 20216 34345 20244
rect 34112 20204 34118 20216
rect 34333 20213 34345 20216
rect 34379 20213 34391 20247
rect 35710 20244 35716 20256
rect 35671 20216 35716 20244
rect 34333 20207 34391 20213
rect 35710 20204 35716 20216
rect 35768 20204 35774 20256
rect 1104 20154 37628 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 37628 20154
rect 1104 20080 37628 20102
rect 9861 20043 9919 20049
rect 9861 20009 9873 20043
rect 9907 20040 9919 20043
rect 10134 20040 10140 20052
rect 9907 20012 10140 20040
rect 9907 20009 9919 20012
rect 9861 20003 9919 20009
rect 10134 20000 10140 20012
rect 10192 20000 10198 20052
rect 12434 20000 12440 20052
rect 12492 20040 12498 20052
rect 14274 20040 14280 20052
rect 12492 20012 12537 20040
rect 14235 20012 14280 20040
rect 12492 20000 12498 20012
rect 14274 20000 14280 20012
rect 14332 20000 14338 20052
rect 19613 20043 19671 20049
rect 19613 20009 19625 20043
rect 19659 20040 19671 20043
rect 19702 20040 19708 20052
rect 19659 20012 19708 20040
rect 19659 20009 19671 20012
rect 19613 20003 19671 20009
rect 19702 20000 19708 20012
rect 19760 20000 19766 20052
rect 21174 20040 21180 20052
rect 19812 20012 21180 20040
rect 14734 19972 14740 19984
rect 14647 19944 14740 19972
rect 14734 19932 14740 19944
rect 14792 19972 14798 19984
rect 16022 19972 16028 19984
rect 14792 19944 16028 19972
rect 14792 19932 14798 19944
rect 16022 19932 16028 19944
rect 16080 19932 16086 19984
rect 17678 19932 17684 19984
rect 17736 19932 17742 19984
rect 10505 19907 10563 19913
rect 10505 19873 10517 19907
rect 10551 19904 10563 19907
rect 11054 19904 11060 19916
rect 10551 19876 11060 19904
rect 10551 19873 10563 19876
rect 10505 19867 10563 19873
rect 11054 19864 11060 19876
rect 11112 19864 11118 19916
rect 11514 19904 11520 19916
rect 11475 19876 11520 19904
rect 11514 19864 11520 19876
rect 11572 19864 11578 19916
rect 11701 19907 11759 19913
rect 11701 19873 11713 19907
rect 11747 19904 11759 19907
rect 12802 19904 12808 19916
rect 11747 19876 12808 19904
rect 11747 19873 11759 19876
rect 11701 19867 11759 19873
rect 12802 19864 12808 19876
rect 12860 19904 12866 19916
rect 13078 19904 13084 19916
rect 12860 19876 13084 19904
rect 12860 19864 12866 19876
rect 13078 19864 13084 19876
rect 13136 19864 13142 19916
rect 13265 19907 13323 19913
rect 13265 19873 13277 19907
rect 13311 19904 13323 19907
rect 14752 19904 14780 19932
rect 14829 19907 14887 19913
rect 14829 19904 14841 19907
rect 13311 19876 14688 19904
rect 14752 19876 14841 19904
rect 13311 19873 13323 19876
rect 13265 19867 13323 19873
rect 8570 19836 8576 19848
rect 8531 19808 8576 19836
rect 8570 19796 8576 19808
rect 8628 19796 8634 19848
rect 9309 19839 9367 19845
rect 9309 19805 9321 19839
rect 9355 19836 9367 19839
rect 9490 19836 9496 19848
rect 9355 19808 9496 19836
rect 9355 19805 9367 19808
rect 9309 19799 9367 19805
rect 9490 19796 9496 19808
rect 9548 19796 9554 19848
rect 10229 19839 10287 19845
rect 10229 19805 10241 19839
rect 10275 19836 10287 19839
rect 11532 19836 11560 19864
rect 10275 19808 11560 19836
rect 10275 19805 10287 19808
rect 10229 19799 10287 19805
rect 12158 19796 12164 19848
rect 12216 19836 12222 19848
rect 12345 19839 12403 19845
rect 12345 19836 12357 19839
rect 12216 19808 12357 19836
rect 12216 19796 12222 19808
rect 12345 19805 12357 19808
rect 12391 19836 12403 19839
rect 12434 19836 12440 19848
rect 12391 19808 12440 19836
rect 12391 19805 12403 19808
rect 12345 19799 12403 19805
rect 12434 19796 12440 19808
rect 12492 19796 12498 19848
rect 13357 19839 13415 19845
rect 13357 19805 13369 19839
rect 13403 19836 13415 19839
rect 13446 19836 13452 19848
rect 13403 19808 13452 19836
rect 13403 19805 13415 19808
rect 13357 19799 13415 19805
rect 13446 19796 13452 19808
rect 13504 19796 13510 19848
rect 14660 19845 14688 19876
rect 14829 19873 14841 19876
rect 14875 19873 14887 19907
rect 15930 19904 15936 19916
rect 14829 19867 14887 19873
rect 14936 19876 15936 19904
rect 14645 19839 14703 19845
rect 14645 19805 14657 19839
rect 14691 19836 14703 19839
rect 14936 19836 14964 19876
rect 15930 19864 15936 19876
rect 15988 19864 15994 19916
rect 16301 19907 16359 19913
rect 16301 19873 16313 19907
rect 16347 19904 16359 19907
rect 17696 19904 17724 19932
rect 19812 19904 19840 20012
rect 21174 20000 21180 20012
rect 21232 20000 21238 20052
rect 22189 20043 22247 20049
rect 22189 20009 22201 20043
rect 22235 20040 22247 20043
rect 22278 20040 22284 20052
rect 22235 20012 22284 20040
rect 22235 20009 22247 20012
rect 22189 20003 22247 20009
rect 22278 20000 22284 20012
rect 22336 20000 22342 20052
rect 22554 20000 22560 20052
rect 22612 20040 22618 20052
rect 23293 20043 23351 20049
rect 23293 20040 23305 20043
rect 22612 20012 23305 20040
rect 22612 20000 22618 20012
rect 23293 20009 23305 20012
rect 23339 20009 23351 20043
rect 24578 20040 24584 20052
rect 24539 20012 24584 20040
rect 23293 20003 23351 20009
rect 24578 20000 24584 20012
rect 24636 20000 24642 20052
rect 28166 20000 28172 20052
rect 28224 20040 28230 20052
rect 28445 20043 28503 20049
rect 28445 20040 28457 20043
rect 28224 20012 28457 20040
rect 28224 20000 28230 20012
rect 28445 20009 28457 20012
rect 28491 20009 28503 20043
rect 28445 20003 28503 20009
rect 32490 20000 32496 20052
rect 32548 20040 32554 20052
rect 32585 20043 32643 20049
rect 32585 20040 32597 20043
rect 32548 20012 32597 20040
rect 32548 20000 32554 20012
rect 32585 20009 32597 20012
rect 32631 20009 32643 20043
rect 32585 20003 32643 20009
rect 25130 19972 25136 19984
rect 23952 19944 25136 19972
rect 16347 19876 17724 19904
rect 18800 19876 19840 19904
rect 20441 19907 20499 19913
rect 16347 19873 16359 19876
rect 16301 19867 16359 19873
rect 15654 19836 15660 19848
rect 14691 19808 14964 19836
rect 15615 19808 15660 19836
rect 14691 19805 14703 19808
rect 14645 19799 14703 19805
rect 15654 19796 15660 19808
rect 15712 19796 15718 19848
rect 18690 19836 18696 19848
rect 18603 19808 18696 19836
rect 18690 19796 18696 19808
rect 18748 19836 18754 19848
rect 18800 19836 18828 19876
rect 20441 19873 20453 19907
rect 20487 19904 20499 19907
rect 22002 19904 22008 19916
rect 20487 19876 22008 19904
rect 20487 19873 20499 19876
rect 20441 19867 20499 19873
rect 22002 19864 22008 19876
rect 22060 19864 22066 19916
rect 23952 19913 23980 19944
rect 25130 19932 25136 19944
rect 25188 19932 25194 19984
rect 23937 19907 23995 19913
rect 23937 19873 23949 19907
rect 23983 19873 23995 19907
rect 25222 19904 25228 19916
rect 23937 19867 23995 19873
rect 24412 19876 25228 19904
rect 18748 19808 18828 19836
rect 18748 19796 18754 19808
rect 18874 19796 18880 19848
rect 18932 19836 18938 19848
rect 19429 19839 19487 19845
rect 19429 19836 19441 19839
rect 18932 19808 19441 19836
rect 18932 19796 18938 19808
rect 19429 19805 19441 19808
rect 19475 19805 19487 19839
rect 19429 19799 19487 19805
rect 23661 19839 23719 19845
rect 23661 19805 23673 19839
rect 23707 19836 23719 19839
rect 24412 19836 24440 19876
rect 25222 19864 25228 19876
rect 25280 19864 25286 19916
rect 25314 19864 25320 19916
rect 25372 19904 25378 19916
rect 25593 19907 25651 19913
rect 25593 19904 25605 19907
rect 25372 19876 25605 19904
rect 25372 19864 25378 19876
rect 25593 19873 25605 19876
rect 25639 19873 25651 19907
rect 26970 19904 26976 19916
rect 26931 19876 26976 19904
rect 25593 19867 25651 19873
rect 26970 19864 26976 19876
rect 27028 19864 27034 19916
rect 31202 19864 31208 19916
rect 31260 19904 31266 19916
rect 31573 19907 31631 19913
rect 31573 19904 31585 19907
rect 31260 19876 31585 19904
rect 31260 19864 31266 19876
rect 31573 19873 31585 19876
rect 31619 19873 31631 19907
rect 34054 19904 34060 19916
rect 34015 19876 34060 19904
rect 31573 19867 31631 19873
rect 34054 19864 34060 19876
rect 34112 19864 34118 19916
rect 34330 19904 34336 19916
rect 34291 19876 34336 19904
rect 34330 19864 34336 19876
rect 34388 19864 34394 19916
rect 24762 19836 24768 19848
rect 23707 19808 24440 19836
rect 24723 19808 24768 19836
rect 23707 19805 23719 19808
rect 23661 19799 23719 19805
rect 24762 19796 24768 19808
rect 24820 19796 24826 19848
rect 26418 19796 26424 19848
rect 26476 19836 26482 19848
rect 26697 19839 26755 19845
rect 26697 19836 26709 19839
rect 26476 19808 26709 19836
rect 26476 19796 26482 19808
rect 26697 19805 26709 19808
rect 26743 19805 26755 19839
rect 26697 19799 26755 19805
rect 9582 19728 9588 19780
rect 9640 19768 9646 19780
rect 10321 19771 10379 19777
rect 10321 19768 10333 19771
rect 9640 19740 10333 19768
rect 9640 19728 9646 19740
rect 10321 19737 10333 19740
rect 10367 19737 10379 19771
rect 10321 19731 10379 19737
rect 11425 19771 11483 19777
rect 11425 19737 11437 19771
rect 11471 19768 11483 19771
rect 11606 19768 11612 19780
rect 11471 19740 11612 19768
rect 11471 19737 11483 19740
rect 11425 19731 11483 19737
rect 11606 19728 11612 19740
rect 11664 19728 11670 19780
rect 14458 19728 14464 19780
rect 14516 19768 14522 19780
rect 14737 19771 14795 19777
rect 14737 19768 14749 19771
rect 14516 19740 14749 19768
rect 14516 19728 14522 19740
rect 14737 19737 14749 19740
rect 14783 19737 14795 19771
rect 16577 19771 16635 19777
rect 16577 19768 16589 19771
rect 14737 19731 14795 19737
rect 15856 19740 16589 19768
rect 8386 19700 8392 19712
rect 8347 19672 8392 19700
rect 8386 19660 8392 19672
rect 8444 19660 8450 19712
rect 9217 19703 9275 19709
rect 9217 19669 9229 19703
rect 9263 19700 9275 19703
rect 9306 19700 9312 19712
rect 9263 19672 9312 19700
rect 9263 19669 9275 19672
rect 9217 19663 9275 19669
rect 9306 19660 9312 19672
rect 9364 19660 9370 19712
rect 10594 19660 10600 19712
rect 10652 19700 10658 19712
rect 11057 19703 11115 19709
rect 11057 19700 11069 19703
rect 10652 19672 11069 19700
rect 10652 19660 10658 19672
rect 11057 19669 11069 19672
rect 11103 19669 11115 19703
rect 13722 19700 13728 19712
rect 13683 19672 13728 19700
rect 11057 19663 11115 19669
rect 13722 19660 13728 19672
rect 13780 19660 13786 19712
rect 15856 19709 15884 19740
rect 16577 19737 16589 19740
rect 16623 19737 16635 19771
rect 16577 19731 16635 19737
rect 17586 19728 17592 19780
rect 17644 19728 17650 19780
rect 20714 19768 20720 19780
rect 20675 19740 20720 19768
rect 20714 19728 20720 19740
rect 20772 19728 20778 19780
rect 21266 19728 21272 19780
rect 21324 19728 21330 19780
rect 28258 19768 28264 19780
rect 22066 19740 27384 19768
rect 28198 19740 28264 19768
rect 15841 19703 15899 19709
rect 15841 19669 15853 19703
rect 15887 19669 15899 19703
rect 15841 19663 15899 19669
rect 17954 19660 17960 19712
rect 18012 19700 18018 19712
rect 18049 19703 18107 19709
rect 18049 19700 18061 19703
rect 18012 19672 18061 19700
rect 18012 19660 18018 19672
rect 18049 19669 18061 19672
rect 18095 19669 18107 19703
rect 18782 19700 18788 19712
rect 18743 19672 18788 19700
rect 18049 19663 18107 19669
rect 18782 19660 18788 19672
rect 18840 19660 18846 19712
rect 18966 19660 18972 19712
rect 19024 19700 19030 19712
rect 22066 19700 22094 19740
rect 23750 19700 23756 19712
rect 19024 19672 22094 19700
rect 23711 19672 23756 19700
rect 19024 19660 19030 19672
rect 23750 19660 23756 19672
rect 23808 19660 23814 19712
rect 25038 19660 25044 19712
rect 25096 19700 25102 19712
rect 25777 19703 25835 19709
rect 25777 19700 25789 19703
rect 25096 19672 25789 19700
rect 25096 19660 25102 19672
rect 25777 19669 25789 19672
rect 25823 19669 25835 19703
rect 25777 19663 25835 19669
rect 25866 19660 25872 19712
rect 25924 19700 25930 19712
rect 26237 19703 26295 19709
rect 25924 19672 25969 19700
rect 25924 19660 25930 19672
rect 26237 19669 26249 19703
rect 26283 19700 26295 19703
rect 26786 19700 26792 19712
rect 26283 19672 26792 19700
rect 26283 19669 26295 19672
rect 26237 19663 26295 19669
rect 26786 19660 26792 19672
rect 26844 19660 26850 19712
rect 27356 19700 27384 19740
rect 28258 19728 28264 19740
rect 28316 19728 28322 19780
rect 30834 19728 30840 19780
rect 30892 19728 30898 19780
rect 31294 19768 31300 19780
rect 31255 19740 31300 19768
rect 31294 19728 31300 19740
rect 31352 19728 31358 19780
rect 35710 19768 35716 19780
rect 33626 19740 35716 19768
rect 35710 19728 35716 19740
rect 35768 19728 35774 19780
rect 29730 19700 29736 19712
rect 27356 19672 29736 19700
rect 29730 19660 29736 19672
rect 29788 19700 29794 19712
rect 29825 19703 29883 19709
rect 29825 19700 29837 19703
rect 29788 19672 29837 19700
rect 29788 19660 29794 19672
rect 29825 19669 29837 19672
rect 29871 19669 29883 19703
rect 29825 19663 29883 19669
rect 1104 19610 37628 19632
rect 1104 19558 4874 19610
rect 4926 19558 4938 19610
rect 4990 19558 5002 19610
rect 5054 19558 5066 19610
rect 5118 19558 5130 19610
rect 5182 19558 35594 19610
rect 35646 19558 35658 19610
rect 35710 19558 35722 19610
rect 35774 19558 35786 19610
rect 35838 19558 35850 19610
rect 35902 19558 37628 19610
rect 1104 19536 37628 19558
rect 8570 19456 8576 19508
rect 8628 19496 8634 19508
rect 10229 19499 10287 19505
rect 10229 19496 10241 19499
rect 8628 19468 10241 19496
rect 8628 19456 8634 19468
rect 10229 19465 10241 19468
rect 10275 19465 10287 19499
rect 10594 19496 10600 19508
rect 10555 19468 10600 19496
rect 10229 19459 10287 19465
rect 10594 19456 10600 19468
rect 10652 19456 10658 19508
rect 12989 19499 13047 19505
rect 12989 19496 13001 19499
rect 12360 19468 13001 19496
rect 8294 19428 8300 19440
rect 8036 19400 8300 19428
rect 8036 19369 8064 19400
rect 8294 19388 8300 19400
rect 8352 19388 8358 19440
rect 9306 19388 9312 19440
rect 9364 19388 9370 19440
rect 8021 19363 8079 19369
rect 8021 19329 8033 19363
rect 8067 19329 8079 19363
rect 8021 19323 8079 19329
rect 9582 19320 9588 19372
rect 9640 19360 9646 19372
rect 10689 19363 10747 19369
rect 10689 19360 10701 19363
rect 9640 19332 10701 19360
rect 9640 19320 9646 19332
rect 8297 19295 8355 19301
rect 8297 19261 8309 19295
rect 8343 19292 8355 19295
rect 8386 19292 8392 19304
rect 8343 19264 8392 19292
rect 8343 19261 8355 19264
rect 8297 19255 8355 19261
rect 8386 19252 8392 19264
rect 8444 19252 8450 19304
rect 9784 19301 9812 19332
rect 10689 19329 10701 19332
rect 10735 19329 10747 19363
rect 11882 19360 11888 19372
rect 11843 19332 11888 19360
rect 10689 19323 10747 19329
rect 11882 19320 11888 19332
rect 11940 19320 11946 19372
rect 12360 19369 12388 19468
rect 12989 19465 13001 19468
rect 13035 19465 13047 19499
rect 12989 19459 13047 19465
rect 13357 19499 13415 19505
rect 13357 19465 13369 19499
rect 13403 19496 13415 19499
rect 13722 19496 13728 19508
rect 13403 19468 13728 19496
rect 13403 19465 13415 19468
rect 13357 19459 13415 19465
rect 13722 19456 13728 19468
rect 13780 19456 13786 19508
rect 15654 19456 15660 19508
rect 15712 19496 15718 19508
rect 16853 19499 16911 19505
rect 16853 19496 16865 19499
rect 15712 19468 16865 19496
rect 15712 19456 15718 19468
rect 16853 19465 16865 19468
rect 16899 19465 16911 19499
rect 16853 19459 16911 19465
rect 17221 19499 17279 19505
rect 17221 19465 17233 19499
rect 17267 19496 17279 19499
rect 18966 19496 18972 19508
rect 17267 19468 18972 19496
rect 17267 19465 17279 19468
rect 17221 19459 17279 19465
rect 18966 19456 18972 19468
rect 19024 19456 19030 19508
rect 20622 19496 20628 19508
rect 20583 19468 20628 19496
rect 20622 19456 20628 19468
rect 20680 19456 20686 19508
rect 20806 19456 20812 19508
rect 20864 19496 20870 19508
rect 20993 19499 21051 19505
rect 20993 19496 21005 19499
rect 20864 19468 21005 19496
rect 20864 19456 20870 19468
rect 20993 19465 21005 19468
rect 21039 19496 21051 19499
rect 22278 19496 22284 19508
rect 21039 19468 22284 19496
rect 21039 19465 21051 19468
rect 20993 19459 21051 19465
rect 22278 19456 22284 19468
rect 22336 19456 22342 19508
rect 23750 19456 23756 19508
rect 23808 19496 23814 19508
rect 23845 19499 23903 19505
rect 23845 19496 23857 19499
rect 23808 19468 23857 19496
rect 23808 19456 23814 19468
rect 23845 19465 23857 19468
rect 23891 19496 23903 19499
rect 24949 19499 25007 19505
rect 23891 19468 24900 19496
rect 23891 19465 23903 19468
rect 23845 19459 23903 19465
rect 12618 19388 12624 19440
rect 12676 19428 12682 19440
rect 14090 19428 14096 19440
rect 12676 19400 14096 19428
rect 12676 19388 12682 19400
rect 14090 19388 14096 19400
rect 14148 19428 14154 19440
rect 14148 19400 14596 19428
rect 14148 19388 14154 19400
rect 12345 19363 12403 19369
rect 12345 19329 12357 19363
rect 12391 19329 12403 19363
rect 12345 19323 12403 19329
rect 13449 19363 13507 19369
rect 13449 19329 13461 19363
rect 13495 19360 13507 19363
rect 14458 19360 14464 19372
rect 13495 19332 14464 19360
rect 13495 19329 13507 19332
rect 13449 19323 13507 19329
rect 14458 19320 14464 19332
rect 14516 19320 14522 19372
rect 14568 19369 14596 19400
rect 15286 19388 15292 19440
rect 15344 19388 15350 19440
rect 18874 19388 18880 19440
rect 18932 19388 18938 19440
rect 21082 19428 21088 19440
rect 21043 19400 21088 19428
rect 21082 19388 21088 19400
rect 21140 19388 21146 19440
rect 22370 19428 22376 19440
rect 22331 19400 22376 19428
rect 22370 19388 22376 19400
rect 22428 19388 22434 19440
rect 24302 19428 24308 19440
rect 23598 19400 24308 19428
rect 24302 19388 24308 19400
rect 24360 19388 24366 19440
rect 14553 19363 14611 19369
rect 14553 19329 14565 19363
rect 14599 19329 14611 19363
rect 14553 19323 14611 19329
rect 19886 19320 19892 19372
rect 19944 19360 19950 19372
rect 19944 19332 19989 19360
rect 19944 19320 19950 19332
rect 22002 19320 22008 19372
rect 22060 19360 22066 19372
rect 22097 19363 22155 19369
rect 22097 19360 22109 19363
rect 22060 19332 22109 19360
rect 22060 19320 22066 19332
rect 22097 19329 22109 19332
rect 22143 19329 22155 19363
rect 24872 19360 24900 19468
rect 24949 19465 24961 19499
rect 24995 19496 25007 19499
rect 25777 19499 25835 19505
rect 25777 19496 25789 19499
rect 24995 19468 25789 19496
rect 24995 19465 25007 19468
rect 24949 19459 25007 19465
rect 25777 19465 25789 19468
rect 25823 19465 25835 19499
rect 25777 19459 25835 19465
rect 26145 19499 26203 19505
rect 26145 19465 26157 19499
rect 26191 19496 26203 19499
rect 27246 19496 27252 19508
rect 26191 19468 27252 19496
rect 26191 19465 26203 19468
rect 26145 19459 26203 19465
rect 25038 19428 25044 19440
rect 24999 19400 25044 19428
rect 25038 19388 25044 19400
rect 25096 19388 25102 19440
rect 26160 19360 26188 19459
rect 27246 19456 27252 19468
rect 27304 19456 27310 19508
rect 28905 19499 28963 19505
rect 28905 19496 28917 19499
rect 27816 19468 28917 19496
rect 27816 19428 27844 19468
rect 28905 19465 28917 19468
rect 28951 19496 28963 19499
rect 28994 19496 29000 19508
rect 28951 19468 29000 19496
rect 28951 19465 28963 19468
rect 28905 19459 28963 19465
rect 28994 19456 29000 19468
rect 29052 19456 29058 19508
rect 30834 19496 30840 19508
rect 30795 19468 30840 19496
rect 30834 19456 30840 19468
rect 30892 19456 30898 19508
rect 29457 19431 29515 19437
rect 29457 19428 29469 19431
rect 24872 19332 26188 19360
rect 26252 19400 27844 19428
rect 28658 19400 29469 19428
rect 22097 19323 22155 19329
rect 9769 19295 9827 19301
rect 9769 19261 9781 19295
rect 9815 19261 9827 19295
rect 9769 19255 9827 19261
rect 10781 19295 10839 19301
rect 10781 19261 10793 19295
rect 10827 19261 10839 19295
rect 10781 19255 10839 19261
rect 10686 19184 10692 19236
rect 10744 19224 10750 19236
rect 10796 19224 10824 19255
rect 12710 19252 12716 19304
rect 12768 19292 12774 19304
rect 13541 19295 13599 19301
rect 13541 19292 13553 19295
rect 12768 19264 13553 19292
rect 12768 19252 12774 19264
rect 13541 19261 13553 19264
rect 13587 19292 13599 19295
rect 13630 19292 13636 19304
rect 13587 19264 13636 19292
rect 13587 19261 13599 19264
rect 13541 19255 13599 19261
rect 13630 19252 13636 19264
rect 13688 19252 13694 19304
rect 13722 19252 13728 19304
rect 13780 19292 13786 19304
rect 14829 19295 14887 19301
rect 14829 19292 14841 19295
rect 13780 19264 14841 19292
rect 13780 19252 13786 19264
rect 14829 19261 14841 19264
rect 14875 19261 14887 19295
rect 17310 19292 17316 19304
rect 17271 19264 17316 19292
rect 14829 19255 14887 19261
rect 17310 19252 17316 19264
rect 17368 19252 17374 19304
rect 17405 19295 17463 19301
rect 17405 19261 17417 19295
rect 17451 19261 17463 19295
rect 17405 19255 17463 19261
rect 10744 19196 10824 19224
rect 16301 19227 16359 19233
rect 10744 19184 10750 19196
rect 16301 19193 16313 19227
rect 16347 19224 16359 19227
rect 16482 19224 16488 19236
rect 16347 19196 16488 19224
rect 16347 19193 16359 19196
rect 16301 19187 16359 19193
rect 16482 19184 16488 19196
rect 16540 19224 16546 19236
rect 17420 19224 17448 19255
rect 19150 19252 19156 19304
rect 19208 19292 19214 19304
rect 19613 19295 19671 19301
rect 19613 19292 19625 19295
rect 19208 19264 19625 19292
rect 19208 19252 19214 19264
rect 19613 19261 19625 19264
rect 19659 19261 19671 19295
rect 19613 19255 19671 19261
rect 20254 19252 20260 19304
rect 20312 19292 20318 19304
rect 21177 19295 21235 19301
rect 21177 19292 21189 19295
rect 20312 19264 21189 19292
rect 20312 19252 20318 19264
rect 21177 19261 21189 19264
rect 21223 19261 21235 19295
rect 25130 19292 25136 19304
rect 25091 19264 25136 19292
rect 21177 19255 21235 19261
rect 25130 19252 25136 19264
rect 25188 19252 25194 19304
rect 25866 19252 25872 19304
rect 25924 19292 25930 19304
rect 26252 19301 26280 19400
rect 29457 19397 29469 19400
rect 29503 19397 29515 19431
rect 29457 19391 29515 19397
rect 32766 19388 32772 19440
rect 32824 19388 32830 19440
rect 26418 19320 26424 19372
rect 26476 19360 26482 19372
rect 27157 19363 27215 19369
rect 27157 19360 27169 19363
rect 26476 19332 27169 19360
rect 26476 19320 26482 19332
rect 27157 19329 27169 19332
rect 27203 19329 27215 19363
rect 27157 19323 27215 19329
rect 28718 19320 28724 19372
rect 28776 19360 28782 19372
rect 29549 19363 29607 19369
rect 29549 19360 29561 19363
rect 28776 19332 29561 19360
rect 28776 19320 28782 19332
rect 29549 19329 29561 19332
rect 29595 19329 29607 19363
rect 29549 19323 29607 19329
rect 30558 19320 30564 19372
rect 30616 19360 30622 19372
rect 30929 19363 30987 19369
rect 30929 19360 30941 19363
rect 30616 19332 30941 19360
rect 30616 19320 30622 19332
rect 30929 19329 30941 19332
rect 30975 19360 30987 19363
rect 31570 19360 31576 19372
rect 30975 19332 31576 19360
rect 30975 19329 30987 19332
rect 30929 19323 30987 19329
rect 31570 19320 31576 19332
rect 31628 19320 31634 19372
rect 34057 19363 34115 19369
rect 34057 19329 34069 19363
rect 34103 19360 34115 19363
rect 34330 19360 34336 19372
rect 34103 19332 34336 19360
rect 34103 19329 34115 19332
rect 34057 19323 34115 19329
rect 34330 19320 34336 19332
rect 34388 19320 34394 19372
rect 26237 19295 26295 19301
rect 26237 19292 26249 19295
rect 25924 19264 26249 19292
rect 25924 19252 25930 19264
rect 26237 19261 26249 19264
rect 26283 19261 26295 19295
rect 26237 19255 26295 19261
rect 26329 19295 26387 19301
rect 26329 19261 26341 19295
rect 26375 19261 26387 19295
rect 26329 19255 26387 19261
rect 16540 19196 17448 19224
rect 16540 19184 16546 19196
rect 25774 19184 25780 19236
rect 25832 19224 25838 19236
rect 26344 19224 26372 19255
rect 26970 19252 26976 19304
rect 27028 19292 27034 19304
rect 27433 19295 27491 19301
rect 27433 19292 27445 19295
rect 27028 19264 27445 19292
rect 27028 19252 27034 19264
rect 27433 19261 27445 19264
rect 27479 19261 27491 19295
rect 27433 19255 27491 19261
rect 31018 19252 31024 19304
rect 31076 19292 31082 19304
rect 33781 19295 33839 19301
rect 33781 19292 33793 19295
rect 31076 19264 33793 19292
rect 31076 19252 31082 19264
rect 33781 19261 33793 19264
rect 33827 19261 33839 19295
rect 33781 19255 33839 19261
rect 25832 19196 26372 19224
rect 25832 19184 25838 19196
rect 11698 19156 11704 19168
rect 11659 19128 11704 19156
rect 11698 19116 11704 19128
rect 11756 19116 11762 19168
rect 12529 19159 12587 19165
rect 12529 19125 12541 19159
rect 12575 19156 12587 19159
rect 12894 19156 12900 19168
rect 12575 19128 12900 19156
rect 12575 19125 12587 19128
rect 12529 19119 12587 19125
rect 12894 19116 12900 19128
rect 12952 19116 12958 19168
rect 18046 19116 18052 19168
rect 18104 19156 18110 19168
rect 18141 19159 18199 19165
rect 18141 19156 18153 19159
rect 18104 19128 18153 19156
rect 18104 19116 18110 19128
rect 18141 19125 18153 19128
rect 18187 19125 18199 19159
rect 18141 19119 18199 19125
rect 23934 19116 23940 19168
rect 23992 19156 23998 19168
rect 24581 19159 24639 19165
rect 24581 19156 24593 19159
rect 23992 19128 24593 19156
rect 23992 19116 23998 19128
rect 24581 19125 24593 19128
rect 24627 19125 24639 19159
rect 24581 19119 24639 19125
rect 28442 19116 28448 19168
rect 28500 19156 28506 19168
rect 31386 19156 31392 19168
rect 28500 19128 31392 19156
rect 28500 19116 28506 19128
rect 31386 19116 31392 19128
rect 31444 19116 31450 19168
rect 31846 19116 31852 19168
rect 31904 19156 31910 19168
rect 32309 19159 32367 19165
rect 32309 19156 32321 19159
rect 31904 19128 32321 19156
rect 31904 19116 31910 19128
rect 32309 19125 32321 19128
rect 32355 19125 32367 19159
rect 32309 19119 32367 19125
rect 1104 19066 37628 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 37628 19066
rect 1104 18992 37628 19014
rect 1762 18912 1768 18964
rect 1820 18952 1826 18964
rect 7006 18952 7012 18964
rect 1820 18924 7012 18952
rect 1820 18912 1826 18924
rect 7006 18912 7012 18924
rect 7064 18952 7070 18964
rect 7745 18955 7803 18961
rect 7745 18952 7757 18955
rect 7064 18924 7757 18952
rect 7064 18912 7070 18924
rect 7745 18921 7757 18924
rect 7791 18921 7803 18955
rect 7745 18915 7803 18921
rect 11882 18912 11888 18964
rect 11940 18952 11946 18964
rect 12069 18955 12127 18961
rect 12069 18952 12081 18955
rect 11940 18924 12081 18952
rect 11940 18912 11946 18924
rect 12069 18921 12081 18924
rect 12115 18921 12127 18955
rect 13722 18952 13728 18964
rect 13683 18924 13728 18952
rect 12069 18915 12127 18921
rect 13722 18912 13728 18924
rect 13780 18912 13786 18964
rect 14369 18955 14427 18961
rect 14369 18921 14381 18955
rect 14415 18952 14427 18955
rect 15286 18952 15292 18964
rect 14415 18924 15292 18952
rect 14415 18921 14427 18924
rect 14369 18915 14427 18921
rect 15286 18912 15292 18924
rect 15344 18912 15350 18964
rect 15654 18912 15660 18964
rect 15712 18952 15718 18964
rect 17037 18955 17095 18961
rect 17037 18952 17049 18955
rect 15712 18924 17049 18952
rect 15712 18912 15718 18924
rect 17037 18921 17049 18924
rect 17083 18921 17095 18955
rect 17037 18915 17095 18921
rect 18785 18955 18843 18961
rect 18785 18921 18797 18955
rect 18831 18952 18843 18955
rect 18874 18952 18880 18964
rect 18831 18924 18880 18952
rect 18831 18921 18843 18924
rect 18785 18915 18843 18921
rect 18874 18912 18880 18924
rect 18932 18912 18938 18964
rect 19426 18952 19432 18964
rect 19387 18924 19432 18952
rect 19426 18912 19432 18924
rect 19484 18912 19490 18964
rect 25038 18912 25044 18964
rect 25096 18952 25102 18964
rect 26329 18955 26387 18961
rect 26329 18952 26341 18955
rect 25096 18924 26341 18952
rect 25096 18912 25102 18924
rect 26329 18921 26341 18924
rect 26375 18921 26387 18955
rect 26970 18952 26976 18964
rect 26931 18924 26976 18952
rect 26329 18915 26387 18921
rect 26970 18912 26976 18924
rect 27028 18912 27034 18964
rect 31018 18952 31024 18964
rect 30979 18924 31024 18952
rect 31018 18912 31024 18924
rect 31076 18912 31082 18964
rect 32766 18912 32772 18964
rect 32824 18952 32830 18964
rect 32861 18955 32919 18961
rect 32861 18952 32873 18955
rect 32824 18924 32873 18952
rect 32824 18912 32830 18924
rect 32861 18921 32873 18924
rect 32907 18921 32919 18955
rect 32861 18915 32919 18921
rect 16574 18844 16580 18896
rect 16632 18884 16638 18896
rect 19794 18884 19800 18896
rect 16632 18856 19800 18884
rect 16632 18844 16638 18856
rect 19794 18844 19800 18856
rect 19852 18844 19858 18896
rect 29196 18856 30880 18884
rect 5997 18819 6055 18825
rect 5997 18785 6009 18819
rect 6043 18816 6055 18819
rect 8294 18816 8300 18828
rect 6043 18788 8300 18816
rect 6043 18785 6055 18788
rect 5997 18779 6055 18785
rect 8294 18776 8300 18788
rect 8352 18816 8358 18828
rect 9125 18819 9183 18825
rect 9125 18816 9137 18819
rect 8352 18788 9137 18816
rect 8352 18776 8358 18788
rect 9125 18785 9137 18788
rect 9171 18816 9183 18819
rect 9398 18816 9404 18828
rect 9171 18788 9404 18816
rect 9171 18785 9183 18788
rect 9125 18779 9183 18785
rect 9398 18776 9404 18788
rect 9456 18776 9462 18828
rect 11054 18776 11060 18828
rect 11112 18816 11118 18828
rect 11425 18819 11483 18825
rect 11425 18816 11437 18819
rect 11112 18788 11437 18816
rect 11112 18776 11118 18788
rect 11425 18785 11437 18788
rect 11471 18785 11483 18819
rect 11606 18816 11612 18828
rect 11567 18788 11612 18816
rect 11425 18779 11483 18785
rect 11440 18748 11468 18779
rect 11606 18776 11612 18788
rect 11664 18776 11670 18828
rect 12434 18776 12440 18828
rect 12492 18816 12498 18828
rect 13722 18816 13728 18828
rect 12492 18788 13728 18816
rect 12492 18776 12498 18788
rect 12912 18757 12940 18788
rect 13722 18776 13728 18788
rect 13780 18776 13786 18828
rect 15565 18819 15623 18825
rect 15565 18785 15577 18819
rect 15611 18816 15623 18819
rect 16206 18816 16212 18828
rect 15611 18788 16212 18816
rect 15611 18785 15623 18788
rect 15565 18779 15623 18785
rect 16206 18776 16212 18788
rect 16264 18816 16270 18828
rect 16942 18816 16948 18828
rect 16264 18788 16948 18816
rect 16264 18776 16270 18788
rect 16942 18776 16948 18788
rect 17000 18776 17006 18828
rect 17681 18819 17739 18825
rect 17681 18785 17693 18819
rect 17727 18816 17739 18819
rect 20254 18816 20260 18828
rect 17727 18788 20260 18816
rect 17727 18785 17739 18788
rect 17681 18779 17739 18785
rect 12897 18751 12955 18757
rect 11440 18720 12434 18748
rect 5994 18640 6000 18692
rect 6052 18680 6058 18692
rect 6273 18683 6331 18689
rect 6273 18680 6285 18683
rect 6052 18652 6285 18680
rect 6052 18640 6058 18652
rect 6273 18649 6285 18652
rect 6319 18649 6331 18683
rect 6273 18643 6331 18649
rect 7282 18640 7288 18692
rect 7340 18640 7346 18692
rect 8386 18640 8392 18692
rect 8444 18680 8450 18692
rect 9401 18683 9459 18689
rect 9401 18680 9413 18683
rect 8444 18652 9413 18680
rect 8444 18640 8450 18652
rect 9401 18649 9413 18652
rect 9447 18649 9459 18683
rect 9401 18643 9459 18649
rect 9858 18640 9864 18692
rect 9916 18640 9922 18692
rect 12406 18680 12434 18720
rect 12897 18717 12909 18751
rect 12943 18717 12955 18751
rect 13538 18748 13544 18760
rect 13499 18720 13544 18748
rect 12897 18711 12955 18717
rect 13538 18708 13544 18720
rect 13596 18708 13602 18760
rect 14274 18748 14280 18760
rect 14235 18720 14280 18748
rect 14274 18708 14280 18720
rect 14332 18708 14338 18760
rect 14458 18708 14464 18760
rect 14516 18748 14522 18760
rect 15289 18751 15347 18757
rect 15289 18748 15301 18751
rect 14516 18720 15301 18748
rect 14516 18708 14522 18720
rect 15289 18717 15301 18720
rect 15335 18717 15347 18751
rect 15289 18711 15347 18717
rect 15381 18751 15439 18757
rect 15381 18717 15393 18751
rect 15427 18748 15439 18751
rect 16482 18748 16488 18760
rect 15427 18720 16488 18748
rect 15427 18717 15439 18720
rect 15381 18711 15439 18717
rect 16482 18708 16488 18720
rect 16540 18708 16546 18760
rect 17310 18708 17316 18760
rect 17368 18748 17374 18760
rect 17405 18751 17463 18757
rect 17405 18748 17417 18751
rect 17368 18720 17417 18748
rect 17368 18708 17374 18720
rect 17405 18717 17417 18720
rect 17451 18717 17463 18751
rect 17405 18711 17463 18717
rect 13354 18680 13360 18692
rect 12406 18652 13360 18680
rect 13354 18640 13360 18652
rect 13412 18640 13418 18692
rect 15470 18640 15476 18692
rect 15528 18680 15534 18692
rect 17696 18680 17724 18779
rect 20254 18776 20260 18788
rect 20312 18776 20318 18828
rect 21177 18819 21235 18825
rect 21177 18785 21189 18819
rect 21223 18816 21235 18819
rect 22002 18816 22008 18828
rect 21223 18788 22008 18816
rect 21223 18785 21235 18788
rect 21177 18779 21235 18785
rect 22002 18776 22008 18788
rect 22060 18816 22066 18828
rect 24581 18819 24639 18825
rect 24581 18816 24593 18819
rect 22060 18788 24593 18816
rect 22060 18776 22066 18788
rect 24581 18785 24593 18788
rect 24627 18785 24639 18819
rect 24581 18779 24639 18785
rect 29196 18760 29224 18856
rect 30742 18816 30748 18828
rect 29840 18788 30748 18816
rect 17770 18708 17776 18760
rect 17828 18748 17834 18760
rect 18877 18751 18935 18757
rect 18877 18748 18889 18751
rect 17828 18720 18889 18748
rect 17828 18708 17834 18720
rect 18877 18717 18889 18720
rect 18923 18717 18935 18751
rect 18877 18711 18935 18717
rect 22094 18708 22100 18760
rect 22152 18748 22158 18760
rect 22833 18751 22891 18757
rect 22152 18720 22197 18748
rect 22152 18708 22158 18720
rect 22833 18717 22845 18751
rect 22879 18717 22891 18751
rect 22833 18711 22891 18717
rect 23845 18751 23903 18757
rect 23845 18717 23857 18751
rect 23891 18748 23903 18751
rect 23934 18748 23940 18760
rect 23891 18720 23940 18748
rect 23891 18717 23903 18720
rect 23845 18711 23903 18717
rect 15528 18652 17724 18680
rect 15528 18640 15534 18652
rect 18782 18640 18788 18692
rect 18840 18680 18846 18692
rect 20898 18680 20904 18692
rect 18840 18652 19734 18680
rect 20859 18652 20904 18680
rect 18840 18640 18846 18652
rect 20898 18640 20904 18652
rect 20956 18640 20962 18692
rect 21821 18683 21879 18689
rect 21821 18649 21833 18683
rect 21867 18680 21879 18683
rect 21910 18680 21916 18692
rect 21867 18652 21916 18680
rect 21867 18649 21879 18652
rect 21821 18643 21879 18649
rect 21910 18640 21916 18652
rect 21968 18680 21974 18692
rect 22848 18680 22876 18711
rect 23934 18708 23940 18720
rect 23992 18708 23998 18760
rect 26786 18748 26792 18760
rect 26747 18720 26792 18748
rect 26786 18708 26792 18720
rect 26844 18708 26850 18760
rect 27522 18708 27528 18760
rect 27580 18748 27586 18760
rect 27617 18751 27675 18757
rect 27617 18748 27629 18751
rect 27580 18720 27629 18748
rect 27580 18708 27586 18720
rect 27617 18717 27629 18720
rect 27663 18717 27675 18751
rect 28994 18748 29000 18760
rect 28955 18720 29000 18748
rect 27617 18711 27675 18717
rect 28994 18708 29000 18720
rect 29052 18708 29058 18760
rect 29178 18748 29184 18760
rect 29139 18720 29184 18748
rect 29178 18708 29184 18720
rect 29236 18708 29242 18760
rect 29840 18757 29868 18788
rect 30742 18776 30748 18788
rect 30800 18776 30806 18828
rect 29825 18751 29883 18757
rect 29825 18717 29837 18751
rect 29871 18717 29883 18751
rect 29825 18711 29883 18717
rect 30009 18751 30067 18757
rect 30009 18717 30021 18751
rect 30055 18717 30067 18751
rect 30009 18711 30067 18717
rect 30653 18751 30711 18757
rect 30653 18717 30665 18751
rect 30699 18748 30711 18751
rect 30852 18748 30880 18856
rect 32125 18819 32183 18825
rect 32125 18785 32137 18819
rect 32171 18816 32183 18819
rect 32171 18788 32812 18816
rect 32171 18785 32183 18788
rect 32125 18779 32183 18785
rect 31846 18748 31852 18760
rect 30699 18720 31852 18748
rect 30699 18717 30711 18720
rect 30653 18711 30711 18717
rect 24857 18683 24915 18689
rect 24857 18680 24869 18683
rect 21968 18652 22876 18680
rect 24044 18652 24869 18680
rect 21968 18640 21974 18652
rect 2038 18572 2044 18624
rect 2096 18612 2102 18624
rect 9674 18612 9680 18624
rect 2096 18584 9680 18612
rect 2096 18572 2102 18584
rect 9674 18572 9680 18584
rect 9732 18612 9738 18624
rect 10873 18615 10931 18621
rect 10873 18612 10885 18615
rect 9732 18584 10885 18612
rect 9732 18572 9738 18584
rect 10873 18581 10885 18584
rect 10919 18581 10931 18615
rect 10873 18575 10931 18581
rect 11701 18615 11759 18621
rect 11701 18581 11713 18615
rect 11747 18612 11759 18615
rect 12158 18612 12164 18624
rect 11747 18584 12164 18612
rect 11747 18581 11759 18584
rect 11701 18575 11759 18581
rect 12158 18572 12164 18584
rect 12216 18572 12222 18624
rect 12986 18612 12992 18624
rect 12947 18584 12992 18612
rect 12986 18572 12992 18584
rect 13044 18572 13050 18624
rect 14918 18612 14924 18624
rect 14879 18584 14924 18612
rect 14918 18572 14924 18584
rect 14976 18572 14982 18624
rect 15194 18572 15200 18624
rect 15252 18612 15258 18624
rect 16209 18615 16267 18621
rect 16209 18612 16221 18615
rect 15252 18584 16221 18612
rect 15252 18572 15258 18584
rect 16209 18581 16221 18584
rect 16255 18612 16267 18615
rect 16574 18612 16580 18624
rect 16255 18584 16580 18612
rect 16255 18581 16267 18584
rect 16209 18575 16267 18581
rect 16574 18572 16580 18584
rect 16632 18572 16638 18624
rect 17494 18572 17500 18624
rect 17552 18612 17558 18624
rect 22922 18612 22928 18624
rect 17552 18584 17597 18612
rect 22883 18584 22928 18612
rect 17552 18572 17558 18584
rect 22922 18572 22928 18584
rect 22980 18572 22986 18624
rect 24044 18621 24072 18652
rect 24857 18649 24869 18652
rect 24903 18649 24915 18683
rect 24857 18643 24915 18649
rect 25314 18640 25320 18692
rect 25372 18640 25378 18692
rect 28350 18680 28356 18692
rect 28311 18652 28356 18680
rect 28350 18640 28356 18652
rect 28408 18640 28414 18692
rect 30024 18680 30052 18711
rect 31846 18708 31852 18720
rect 31904 18708 31910 18760
rect 32306 18748 32312 18760
rect 32267 18720 32312 18748
rect 32306 18708 32312 18720
rect 32364 18708 32370 18760
rect 32784 18757 32812 18788
rect 32769 18751 32827 18757
rect 32769 18717 32781 18751
rect 32815 18748 32827 18751
rect 33410 18748 33416 18760
rect 32815 18720 33416 18748
rect 32815 18717 32827 18720
rect 32769 18711 32827 18717
rect 33410 18708 33416 18720
rect 33468 18748 33474 18760
rect 35069 18751 35127 18757
rect 35069 18748 35081 18751
rect 33468 18720 35081 18748
rect 33468 18708 33474 18720
rect 35069 18717 35081 18720
rect 35115 18717 35127 18751
rect 35069 18711 35127 18717
rect 31294 18680 31300 18692
rect 30024 18652 31300 18680
rect 31294 18640 31300 18652
rect 31352 18640 31358 18692
rect 24029 18615 24087 18621
rect 24029 18581 24041 18615
rect 24075 18581 24087 18615
rect 24029 18575 24087 18581
rect 28810 18572 28816 18624
rect 28868 18612 28874 18624
rect 28997 18615 29055 18621
rect 28997 18612 29009 18615
rect 28868 18584 29009 18612
rect 28868 18572 28874 18584
rect 28997 18581 29009 18584
rect 29043 18581 29055 18615
rect 28997 18575 29055 18581
rect 29917 18615 29975 18621
rect 29917 18581 29929 18615
rect 29963 18612 29975 18615
rect 30282 18612 30288 18624
rect 29963 18584 30288 18612
rect 29963 18581 29975 18584
rect 29917 18575 29975 18581
rect 30282 18572 30288 18584
rect 30340 18572 30346 18624
rect 34977 18615 35035 18621
rect 34977 18581 34989 18615
rect 35023 18612 35035 18615
rect 35066 18612 35072 18624
rect 35023 18584 35072 18612
rect 35023 18581 35035 18584
rect 34977 18575 35035 18581
rect 35066 18572 35072 18584
rect 35124 18572 35130 18624
rect 1104 18522 37628 18544
rect 1104 18470 4874 18522
rect 4926 18470 4938 18522
rect 4990 18470 5002 18522
rect 5054 18470 5066 18522
rect 5118 18470 5130 18522
rect 5182 18470 35594 18522
rect 35646 18470 35658 18522
rect 35710 18470 35722 18522
rect 35774 18470 35786 18522
rect 35838 18470 35850 18522
rect 35902 18470 37628 18522
rect 1104 18448 37628 18470
rect 5994 18408 6000 18420
rect 5955 18380 6000 18408
rect 5994 18368 6000 18380
rect 6052 18368 6058 18420
rect 7193 18411 7251 18417
rect 7193 18377 7205 18411
rect 7239 18408 7251 18411
rect 7282 18408 7288 18420
rect 7239 18380 7288 18408
rect 7239 18377 7251 18380
rect 7193 18371 7251 18377
rect 7282 18368 7288 18380
rect 7340 18368 7346 18420
rect 8205 18411 8263 18417
rect 8205 18377 8217 18411
rect 8251 18408 8263 18411
rect 9858 18408 9864 18420
rect 8251 18380 9864 18408
rect 8251 18377 8263 18380
rect 8205 18371 8263 18377
rect 9858 18368 9864 18380
rect 9916 18368 9922 18420
rect 11146 18408 11152 18420
rect 9968 18380 11008 18408
rect 11059 18380 11152 18408
rect 9766 18340 9772 18352
rect 8128 18312 9772 18340
rect 5813 18275 5871 18281
rect 5813 18241 5825 18275
rect 5859 18272 5871 18275
rect 6362 18272 6368 18284
rect 5859 18244 6368 18272
rect 5859 18241 5871 18244
rect 5813 18235 5871 18241
rect 6362 18232 6368 18244
rect 6420 18232 6426 18284
rect 7282 18272 7288 18284
rect 7195 18244 7288 18272
rect 7282 18232 7288 18244
rect 7340 18272 7346 18284
rect 8128 18281 8156 18312
rect 9766 18300 9772 18312
rect 9824 18340 9830 18352
rect 9968 18340 9996 18380
rect 9824 18312 9996 18340
rect 9824 18300 9830 18312
rect 10134 18300 10140 18352
rect 10192 18300 10198 18352
rect 10980 18340 11008 18380
rect 11146 18368 11152 18380
rect 11204 18408 11210 18420
rect 11606 18408 11612 18420
rect 11204 18380 11612 18408
rect 11204 18368 11210 18380
rect 11606 18368 11612 18380
rect 11664 18368 11670 18420
rect 13538 18368 13544 18420
rect 13596 18408 13602 18420
rect 14829 18411 14887 18417
rect 14829 18408 14841 18411
rect 13596 18380 14841 18408
rect 13596 18368 13602 18380
rect 14829 18377 14841 18380
rect 14875 18377 14887 18411
rect 15194 18408 15200 18420
rect 15155 18380 15200 18408
rect 14829 18371 14887 18377
rect 15194 18368 15200 18380
rect 15252 18368 15258 18420
rect 19061 18411 19119 18417
rect 19061 18408 19073 18411
rect 16132 18380 19073 18408
rect 12894 18340 12900 18352
rect 10980 18312 12020 18340
rect 12855 18312 12900 18340
rect 8113 18275 8171 18281
rect 8113 18272 8125 18275
rect 7340 18244 8125 18272
rect 7340 18232 7346 18244
rect 8113 18241 8125 18244
rect 8159 18241 8171 18275
rect 8113 18235 8171 18241
rect 8757 18275 8815 18281
rect 8757 18241 8769 18275
rect 8803 18272 8815 18275
rect 9214 18272 9220 18284
rect 8803 18244 9220 18272
rect 8803 18241 8815 18244
rect 8757 18235 8815 18241
rect 9214 18232 9220 18244
rect 9272 18232 9278 18284
rect 9398 18272 9404 18284
rect 9359 18244 9404 18272
rect 9398 18232 9404 18244
rect 9456 18232 9462 18284
rect 11992 18281 12020 18312
rect 12894 18300 12900 18312
rect 12952 18300 12958 18352
rect 12986 18300 12992 18352
rect 13044 18340 13050 18352
rect 13044 18312 13386 18340
rect 13044 18300 13050 18312
rect 16132 18281 16160 18380
rect 19061 18377 19073 18380
rect 19107 18377 19119 18411
rect 19426 18408 19432 18420
rect 19387 18380 19432 18408
rect 19061 18371 19119 18377
rect 19426 18368 19432 18380
rect 19484 18368 19490 18420
rect 20806 18408 20812 18420
rect 20767 18380 20812 18408
rect 20806 18368 20812 18380
rect 20864 18368 20870 18420
rect 21910 18368 21916 18420
rect 21968 18408 21974 18420
rect 24305 18411 24363 18417
rect 21968 18380 24256 18408
rect 21968 18368 21974 18380
rect 16574 18300 16580 18352
rect 16632 18340 16638 18352
rect 17129 18343 17187 18349
rect 17129 18340 17141 18343
rect 16632 18312 17141 18340
rect 16632 18300 16638 18312
rect 17129 18309 17141 18312
rect 17175 18309 17187 18343
rect 17129 18303 17187 18309
rect 18138 18300 18144 18352
rect 18196 18300 18202 18352
rect 20898 18340 20904 18352
rect 18616 18312 20904 18340
rect 11977 18275 12035 18281
rect 11977 18241 11989 18275
rect 12023 18241 12035 18275
rect 11977 18235 12035 18241
rect 16117 18275 16175 18281
rect 16117 18241 16129 18275
rect 16163 18241 16175 18275
rect 16117 18235 16175 18241
rect 9677 18207 9735 18213
rect 9677 18204 9689 18207
rect 8956 18176 9689 18204
rect 8956 18145 8984 18176
rect 9677 18173 9689 18176
rect 9723 18173 9735 18207
rect 12618 18204 12624 18216
rect 12579 18176 12624 18204
rect 9677 18167 9735 18173
rect 12618 18164 12624 18176
rect 12676 18164 12682 18216
rect 14369 18207 14427 18213
rect 14369 18173 14381 18207
rect 14415 18204 14427 18207
rect 14458 18204 14464 18216
rect 14415 18176 14464 18204
rect 14415 18173 14427 18176
rect 14369 18167 14427 18173
rect 14458 18164 14464 18176
rect 14516 18164 14522 18216
rect 15286 18204 15292 18216
rect 15247 18176 15292 18204
rect 15286 18164 15292 18176
rect 15344 18164 15350 18216
rect 15470 18204 15476 18216
rect 15431 18176 15476 18204
rect 15470 18164 15476 18176
rect 15528 18164 15534 18216
rect 16758 18164 16764 18216
rect 16816 18204 16822 18216
rect 16853 18207 16911 18213
rect 16853 18204 16865 18207
rect 16816 18176 16865 18204
rect 16816 18164 16822 18176
rect 16853 18173 16865 18176
rect 16899 18173 16911 18207
rect 18616 18204 18644 18312
rect 20898 18300 20904 18312
rect 20956 18300 20962 18352
rect 22922 18300 22928 18352
rect 22980 18300 22986 18352
rect 19521 18275 19579 18281
rect 19521 18241 19533 18275
rect 19567 18272 19579 18275
rect 20714 18272 20720 18284
rect 19567 18244 20720 18272
rect 19567 18241 19579 18244
rect 19521 18235 19579 18241
rect 20714 18232 20720 18244
rect 20772 18232 20778 18284
rect 24228 18281 24256 18380
rect 24305 18377 24317 18411
rect 24351 18408 24363 18411
rect 25314 18408 25320 18420
rect 24351 18380 25320 18408
rect 24351 18377 24363 18380
rect 24305 18371 24363 18377
rect 25314 18368 25320 18380
rect 25372 18368 25378 18420
rect 29454 18408 29460 18420
rect 27172 18380 29460 18408
rect 25038 18300 25044 18352
rect 25096 18340 25102 18352
rect 25225 18343 25283 18349
rect 25225 18340 25237 18343
rect 25096 18312 25237 18340
rect 25096 18300 25102 18312
rect 25225 18309 25237 18312
rect 25271 18309 25283 18343
rect 25225 18303 25283 18309
rect 24213 18275 24271 18281
rect 24213 18241 24225 18275
rect 24259 18241 24271 18275
rect 26050 18272 26056 18284
rect 26011 18244 26056 18272
rect 24213 18235 24271 18241
rect 26050 18232 26056 18244
rect 26108 18232 26114 18284
rect 26786 18232 26792 18284
rect 26844 18272 26850 18284
rect 27172 18281 27200 18380
rect 29454 18368 29460 18380
rect 29512 18368 29518 18420
rect 31202 18408 31208 18420
rect 30116 18380 31208 18408
rect 27433 18343 27491 18349
rect 27433 18309 27445 18343
rect 27479 18340 27491 18343
rect 27522 18340 27528 18352
rect 27479 18312 27528 18340
rect 27479 18309 27491 18312
rect 27433 18303 27491 18309
rect 27157 18275 27215 18281
rect 27157 18272 27169 18275
rect 26844 18244 27169 18272
rect 26844 18232 26850 18244
rect 27157 18241 27169 18244
rect 27203 18241 27215 18275
rect 27157 18235 27215 18241
rect 16853 18167 16911 18173
rect 16960 18176 18644 18204
rect 19705 18207 19763 18213
rect 8941 18139 8999 18145
rect 8941 18105 8953 18139
rect 8987 18105 8999 18139
rect 8941 18099 8999 18105
rect 16301 18139 16359 18145
rect 16301 18105 16313 18139
rect 16347 18136 16359 18139
rect 16960 18136 16988 18176
rect 19705 18173 19717 18207
rect 19751 18204 19763 18207
rect 20254 18204 20260 18216
rect 19751 18176 20260 18204
rect 19751 18173 19763 18176
rect 19705 18167 19763 18173
rect 20254 18164 20260 18176
rect 20312 18164 20318 18216
rect 20990 18204 20996 18216
rect 20951 18176 20996 18204
rect 20990 18164 20996 18176
rect 21048 18164 21054 18216
rect 22002 18204 22008 18216
rect 21963 18176 22008 18204
rect 22002 18164 22008 18176
rect 22060 18164 22066 18216
rect 22278 18204 22284 18216
rect 22239 18176 22284 18204
rect 22278 18164 22284 18176
rect 22336 18164 22342 18216
rect 25314 18204 25320 18216
rect 25275 18176 25320 18204
rect 25314 18164 25320 18176
rect 25372 18164 25378 18216
rect 25498 18164 25504 18216
rect 25556 18204 25562 18216
rect 25774 18204 25780 18216
rect 25556 18176 25780 18204
rect 25556 18164 25562 18176
rect 25774 18164 25780 18176
rect 25832 18164 25838 18216
rect 26970 18164 26976 18216
rect 27028 18204 27034 18216
rect 27448 18204 27476 18303
rect 27522 18300 27528 18312
rect 27580 18300 27586 18352
rect 28810 18340 28816 18352
rect 28771 18312 28816 18340
rect 28810 18300 28816 18312
rect 28868 18300 28874 18352
rect 30116 18340 30144 18380
rect 31202 18368 31208 18380
rect 31260 18368 31266 18420
rect 31754 18368 31760 18420
rect 31812 18408 31818 18420
rect 31812 18380 32352 18408
rect 31812 18368 31818 18380
rect 30282 18340 30288 18352
rect 30024 18312 30144 18340
rect 30243 18312 30288 18340
rect 28534 18272 28540 18284
rect 28495 18244 28540 18272
rect 28534 18232 28540 18244
rect 28592 18232 28598 18284
rect 28626 18232 28632 18284
rect 28684 18272 28690 18284
rect 29086 18281 29092 18284
rect 28905 18275 28963 18281
rect 28684 18244 28729 18272
rect 28684 18232 28690 18244
rect 28905 18241 28917 18275
rect 28951 18241 28963 18275
rect 28905 18235 28963 18241
rect 29043 18275 29092 18281
rect 29043 18241 29055 18275
rect 29089 18241 29092 18275
rect 29043 18235 29092 18241
rect 27028 18176 27476 18204
rect 27028 18164 27034 18176
rect 28074 18164 28080 18216
rect 28132 18204 28138 18216
rect 28920 18204 28948 18235
rect 29086 18232 29092 18235
rect 29144 18232 29150 18284
rect 30024 18281 30052 18312
rect 30282 18300 30288 18312
rect 30340 18300 30346 18352
rect 32324 18349 32352 18380
rect 32398 18368 32404 18420
rect 32456 18408 32462 18420
rect 32493 18411 32551 18417
rect 32493 18408 32505 18411
rect 32456 18380 32505 18408
rect 32456 18368 32462 18380
rect 32493 18377 32505 18380
rect 32539 18377 32551 18411
rect 32493 18371 32551 18377
rect 32309 18343 32367 18349
rect 31510 18312 32260 18340
rect 30009 18275 30067 18281
rect 30009 18241 30021 18275
rect 30055 18241 30067 18275
rect 32232 18272 32260 18312
rect 32309 18309 32321 18343
rect 32355 18309 32367 18343
rect 33137 18343 33195 18349
rect 33137 18340 33149 18343
rect 32309 18303 32367 18309
rect 32416 18312 33149 18340
rect 32416 18272 32444 18312
rect 33137 18309 33149 18312
rect 33183 18309 33195 18343
rect 34330 18340 34336 18352
rect 33137 18303 33195 18309
rect 33796 18312 34336 18340
rect 32232 18244 32444 18272
rect 32585 18275 32643 18281
rect 30009 18235 30067 18241
rect 32585 18241 32597 18275
rect 32631 18241 32643 18275
rect 32585 18235 32643 18241
rect 33229 18275 33287 18281
rect 33229 18241 33241 18275
rect 33275 18272 33287 18275
rect 33410 18272 33416 18284
rect 33275 18244 33416 18272
rect 33275 18241 33287 18244
rect 33229 18235 33287 18241
rect 28132 18176 28948 18204
rect 28132 18164 28138 18176
rect 30374 18164 30380 18216
rect 30432 18204 30438 18216
rect 32600 18204 32628 18235
rect 33410 18232 33416 18244
rect 33468 18232 33474 18284
rect 33796 18281 33824 18312
rect 34330 18300 34336 18312
rect 34388 18300 34394 18352
rect 35066 18300 35072 18352
rect 35124 18300 35130 18352
rect 33781 18275 33839 18281
rect 33781 18241 33793 18275
rect 33827 18241 33839 18275
rect 33781 18235 33839 18241
rect 34054 18204 34060 18216
rect 30432 18176 32628 18204
rect 34015 18176 34060 18204
rect 30432 18164 30438 18176
rect 34054 18164 34060 18176
rect 34112 18164 34118 18216
rect 16347 18108 16988 18136
rect 16347 18105 16359 18108
rect 16301 18099 16359 18105
rect 31294 18096 31300 18148
rect 31352 18136 31358 18148
rect 32309 18139 32367 18145
rect 32309 18136 32321 18139
rect 31352 18108 32321 18136
rect 31352 18096 31358 18108
rect 32309 18105 32321 18108
rect 32355 18105 32367 18139
rect 32309 18099 32367 18105
rect 12066 18068 12072 18080
rect 12027 18040 12072 18068
rect 12066 18028 12072 18040
rect 12124 18028 12130 18080
rect 17310 18028 17316 18080
rect 17368 18068 17374 18080
rect 18601 18071 18659 18077
rect 18601 18068 18613 18071
rect 17368 18040 18613 18068
rect 17368 18028 17374 18040
rect 18601 18037 18613 18040
rect 18647 18037 18659 18071
rect 20346 18068 20352 18080
rect 20307 18040 20352 18068
rect 18601 18031 18659 18037
rect 20346 18028 20352 18040
rect 20404 18028 20410 18080
rect 23658 18028 23664 18080
rect 23716 18068 23722 18080
rect 23753 18071 23811 18077
rect 23753 18068 23765 18071
rect 23716 18040 23765 18068
rect 23716 18028 23722 18040
rect 23753 18037 23765 18040
rect 23799 18037 23811 18071
rect 24854 18068 24860 18080
rect 24815 18040 24860 18068
rect 23753 18031 23811 18037
rect 24854 18028 24860 18040
rect 24912 18028 24918 18080
rect 26237 18071 26295 18077
rect 26237 18037 26249 18071
rect 26283 18068 26295 18071
rect 26694 18068 26700 18080
rect 26283 18040 26700 18068
rect 26283 18037 26295 18040
rect 26237 18031 26295 18037
rect 26694 18028 26700 18040
rect 26752 18028 26758 18080
rect 29181 18071 29239 18077
rect 29181 18037 29193 18071
rect 29227 18068 29239 18071
rect 29454 18068 29460 18080
rect 29227 18040 29460 18068
rect 29227 18037 29239 18040
rect 29181 18031 29239 18037
rect 29454 18028 29460 18040
rect 29512 18028 29518 18080
rect 30926 18028 30932 18080
rect 30984 18068 30990 18080
rect 31754 18068 31760 18080
rect 30984 18040 31760 18068
rect 30984 18028 30990 18040
rect 31754 18028 31760 18040
rect 31812 18028 31818 18080
rect 34790 18028 34796 18080
rect 34848 18068 34854 18080
rect 35529 18071 35587 18077
rect 35529 18068 35541 18071
rect 34848 18040 35541 18068
rect 34848 18028 34854 18040
rect 35529 18037 35541 18040
rect 35575 18037 35587 18071
rect 35529 18031 35587 18037
rect 1104 17978 37628 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 37628 17978
rect 1104 17904 37628 17926
rect 8205 17867 8263 17873
rect 8205 17833 8217 17867
rect 8251 17864 8263 17867
rect 8386 17864 8392 17876
rect 8251 17836 8392 17864
rect 8251 17833 8263 17836
rect 8205 17827 8263 17833
rect 8386 17824 8392 17836
rect 8444 17824 8450 17876
rect 9585 17867 9643 17873
rect 9585 17833 9597 17867
rect 9631 17864 9643 17867
rect 10134 17864 10140 17876
rect 9631 17836 10140 17864
rect 9631 17833 9643 17836
rect 9585 17827 9643 17833
rect 10134 17824 10140 17836
rect 10192 17824 10198 17876
rect 12158 17824 12164 17876
rect 12216 17864 12222 17876
rect 13081 17867 13139 17873
rect 13081 17864 13093 17867
rect 12216 17836 13093 17864
rect 12216 17824 12222 17836
rect 13081 17833 13093 17836
rect 13127 17864 13139 17867
rect 18046 17864 18052 17876
rect 13127 17836 18052 17864
rect 13127 17833 13139 17836
rect 13081 17827 13139 17833
rect 18046 17824 18052 17836
rect 18104 17824 18110 17876
rect 22278 17824 22284 17876
rect 22336 17864 22342 17876
rect 22557 17867 22615 17873
rect 22557 17864 22569 17867
rect 22336 17836 22569 17864
rect 22336 17824 22342 17836
rect 22557 17833 22569 17836
rect 22603 17833 22615 17867
rect 22557 17827 22615 17833
rect 25961 17867 26019 17873
rect 25961 17833 25973 17867
rect 26007 17864 26019 17867
rect 26050 17864 26056 17876
rect 26007 17836 26056 17864
rect 26007 17833 26019 17836
rect 25961 17827 26019 17833
rect 26050 17824 26056 17836
rect 26108 17824 26114 17876
rect 28626 17864 28632 17876
rect 28587 17836 28632 17864
rect 28626 17824 28632 17836
rect 28684 17824 28690 17876
rect 33965 17867 34023 17873
rect 33965 17833 33977 17867
rect 34011 17864 34023 17867
rect 34054 17864 34060 17876
rect 34011 17836 34060 17864
rect 34011 17833 34023 17836
rect 33965 17827 34023 17833
rect 34054 17824 34060 17836
rect 34112 17824 34118 17876
rect 6457 17799 6515 17805
rect 6457 17765 6469 17799
rect 6503 17765 6515 17799
rect 6457 17759 6515 17765
rect 5813 17663 5871 17669
rect 5813 17629 5825 17663
rect 5859 17660 5871 17663
rect 6472 17660 6500 17759
rect 13354 17756 13360 17808
rect 13412 17796 13418 17808
rect 16022 17796 16028 17808
rect 13412 17768 16028 17796
rect 13412 17756 13418 17768
rect 16022 17756 16028 17768
rect 16080 17756 16086 17808
rect 20717 17799 20775 17805
rect 16960 17768 18276 17796
rect 16960 17740 16988 17768
rect 7098 17728 7104 17740
rect 7059 17700 7104 17728
rect 7098 17688 7104 17700
rect 7156 17688 7162 17740
rect 10686 17728 10692 17740
rect 10647 17700 10692 17728
rect 10686 17688 10692 17700
rect 10744 17688 10750 17740
rect 11333 17731 11391 17737
rect 11333 17697 11345 17731
rect 11379 17728 11391 17731
rect 12618 17728 12624 17740
rect 11379 17700 12624 17728
rect 11379 17697 11391 17700
rect 11333 17691 11391 17697
rect 12618 17688 12624 17700
rect 12676 17688 12682 17740
rect 13630 17688 13636 17740
rect 13688 17728 13694 17740
rect 14829 17731 14887 17737
rect 14829 17728 14841 17731
rect 13688 17700 14841 17728
rect 13688 17688 13694 17700
rect 14829 17697 14841 17700
rect 14875 17697 14887 17731
rect 14829 17691 14887 17697
rect 15013 17731 15071 17737
rect 15013 17697 15025 17731
rect 15059 17728 15071 17731
rect 15286 17728 15292 17740
rect 15059 17700 15292 17728
rect 15059 17697 15071 17700
rect 15013 17691 15071 17697
rect 15286 17688 15292 17700
rect 15344 17688 15350 17740
rect 16942 17728 16948 17740
rect 16903 17700 16948 17728
rect 16942 17688 16948 17700
rect 17000 17688 17006 17740
rect 17129 17731 17187 17737
rect 17129 17697 17141 17731
rect 17175 17728 17187 17731
rect 17310 17728 17316 17740
rect 17175 17700 17316 17728
rect 17175 17697 17187 17700
rect 17129 17691 17187 17697
rect 17310 17688 17316 17700
rect 17368 17688 17374 17740
rect 18248 17737 18276 17768
rect 20717 17765 20729 17799
rect 20763 17765 20775 17799
rect 35161 17799 35219 17805
rect 20717 17759 20775 17765
rect 23676 17768 25544 17796
rect 18233 17731 18291 17737
rect 18233 17697 18245 17731
rect 18279 17697 18291 17731
rect 18233 17691 18291 17697
rect 18417 17731 18475 17737
rect 18417 17697 18429 17731
rect 18463 17728 18475 17731
rect 19426 17728 19432 17740
rect 18463 17700 19432 17728
rect 18463 17697 18475 17700
rect 18417 17691 18475 17697
rect 19426 17688 19432 17700
rect 19484 17688 19490 17740
rect 20073 17731 20131 17737
rect 20073 17697 20085 17731
rect 20119 17697 20131 17731
rect 20073 17691 20131 17697
rect 8021 17663 8079 17669
rect 5859 17632 6500 17660
rect 6564 17632 7972 17660
rect 5859 17629 5871 17632
rect 5813 17623 5871 17629
rect 6086 17552 6092 17604
rect 6144 17592 6150 17604
rect 6564 17592 6592 17632
rect 6144 17564 6592 17592
rect 6144 17552 6150 17564
rect 6638 17552 6644 17604
rect 6696 17592 6702 17604
rect 6825 17595 6883 17601
rect 6825 17592 6837 17595
rect 6696 17564 6837 17592
rect 6696 17552 6702 17564
rect 6825 17561 6837 17564
rect 6871 17561 6883 17595
rect 7944 17592 7972 17632
rect 8021 17629 8033 17663
rect 8067 17660 8079 17663
rect 8754 17660 8760 17672
rect 8067 17632 8760 17660
rect 8067 17629 8079 17632
rect 8021 17623 8079 17629
rect 8754 17620 8760 17632
rect 8812 17620 8818 17672
rect 9490 17660 9496 17672
rect 9403 17632 9496 17660
rect 9490 17620 9496 17632
rect 9548 17620 9554 17672
rect 10597 17663 10655 17669
rect 10597 17629 10609 17663
rect 10643 17660 10655 17663
rect 11146 17660 11152 17672
rect 10643 17632 11152 17660
rect 10643 17629 10655 17632
rect 10597 17623 10655 17629
rect 11146 17620 11152 17632
rect 11204 17620 11210 17672
rect 14918 17620 14924 17672
rect 14976 17660 14982 17672
rect 15105 17663 15163 17669
rect 15105 17660 15117 17663
rect 14976 17632 15117 17660
rect 14976 17620 14982 17632
rect 15105 17629 15117 17632
rect 15151 17629 15163 17663
rect 15105 17623 15163 17629
rect 18690 17620 18696 17672
rect 18748 17660 18754 17672
rect 20088 17660 20116 17691
rect 20346 17660 20352 17672
rect 18748 17632 20116 17660
rect 20307 17632 20352 17660
rect 18748 17620 18754 17632
rect 20346 17620 20352 17632
rect 20404 17620 20410 17672
rect 20732 17660 20760 17759
rect 23676 17740 23704 17768
rect 23658 17728 23664 17740
rect 23619 17700 23664 17728
rect 23658 17688 23664 17700
rect 23716 17688 23722 17740
rect 23845 17731 23903 17737
rect 23845 17697 23857 17731
rect 23891 17728 23903 17731
rect 25130 17728 25136 17740
rect 23891 17700 25136 17728
rect 23891 17697 23903 17700
rect 23845 17691 23903 17697
rect 21361 17663 21419 17669
rect 21361 17660 21373 17663
rect 20732 17632 21373 17660
rect 21361 17629 21373 17632
rect 21407 17629 21419 17663
rect 21910 17660 21916 17672
rect 21871 17632 21916 17660
rect 21361 17623 21419 17629
rect 21910 17620 21916 17632
rect 21968 17620 21974 17672
rect 22741 17663 22799 17669
rect 22741 17629 22753 17663
rect 22787 17660 22799 17663
rect 22787 17632 23244 17660
rect 22787 17629 22799 17632
rect 22741 17623 22799 17629
rect 9508 17592 9536 17620
rect 10778 17592 10784 17604
rect 7944 17564 10784 17592
rect 6825 17555 6883 17561
rect 10778 17552 10784 17564
rect 10836 17552 10842 17604
rect 11609 17595 11667 17601
rect 11609 17561 11621 17595
rect 11655 17592 11667 17595
rect 11698 17592 11704 17604
rect 11655 17564 11704 17592
rect 11655 17561 11667 17564
rect 11609 17555 11667 17561
rect 11698 17552 11704 17564
rect 11756 17552 11762 17604
rect 12066 17552 12072 17604
rect 12124 17552 12130 17604
rect 16298 17592 16304 17604
rect 16259 17564 16304 17592
rect 16298 17552 16304 17564
rect 16356 17592 16362 17604
rect 17126 17592 17132 17604
rect 16356 17564 17132 17592
rect 16356 17552 16362 17564
rect 17126 17552 17132 17564
rect 17184 17552 17190 17604
rect 17494 17552 17500 17604
rect 17552 17592 17558 17604
rect 18509 17595 18567 17601
rect 18509 17592 18521 17595
rect 17552 17564 18521 17592
rect 17552 17552 17558 17564
rect 18509 17561 18521 17564
rect 18555 17592 18567 17595
rect 18598 17592 18604 17604
rect 18555 17564 18604 17592
rect 18555 17561 18567 17564
rect 18509 17555 18567 17561
rect 18598 17552 18604 17564
rect 18656 17552 18662 17604
rect 20257 17595 20315 17601
rect 20257 17561 20269 17595
rect 20303 17592 20315 17595
rect 21082 17592 21088 17604
rect 20303 17564 21088 17592
rect 20303 17561 20315 17564
rect 20257 17555 20315 17561
rect 21082 17552 21088 17564
rect 21140 17552 21146 17604
rect 5997 17527 6055 17533
rect 5997 17493 6009 17527
rect 6043 17524 6055 17527
rect 6730 17524 6736 17536
rect 6043 17496 6736 17524
rect 6043 17493 6055 17496
rect 5997 17487 6055 17493
rect 6730 17484 6736 17496
rect 6788 17484 6794 17536
rect 6914 17484 6920 17536
rect 6972 17524 6978 17536
rect 6972 17496 7017 17524
rect 6972 17484 6978 17496
rect 9214 17484 9220 17536
rect 9272 17524 9278 17536
rect 10137 17527 10195 17533
rect 10137 17524 10149 17527
rect 9272 17496 10149 17524
rect 9272 17484 9278 17496
rect 10137 17493 10149 17496
rect 10183 17493 10195 17527
rect 10502 17524 10508 17536
rect 10463 17496 10508 17524
rect 10137 17487 10195 17493
rect 10502 17484 10508 17496
rect 10560 17484 10566 17536
rect 15378 17484 15384 17536
rect 15436 17524 15442 17536
rect 15473 17527 15531 17533
rect 15473 17524 15485 17527
rect 15436 17496 15485 17524
rect 15436 17484 15442 17496
rect 15473 17493 15485 17496
rect 15519 17493 15531 17527
rect 15473 17487 15531 17493
rect 16482 17484 16488 17536
rect 16540 17524 16546 17536
rect 17221 17527 17279 17533
rect 17221 17524 17233 17527
rect 16540 17496 17233 17524
rect 16540 17484 16546 17496
rect 17221 17493 17233 17496
rect 17267 17493 17279 17527
rect 17586 17524 17592 17536
rect 17547 17496 17592 17524
rect 17221 17487 17279 17493
rect 17586 17484 17592 17496
rect 17644 17484 17650 17536
rect 18874 17524 18880 17536
rect 18835 17496 18880 17524
rect 18874 17484 18880 17496
rect 18932 17484 18938 17536
rect 21174 17524 21180 17536
rect 21135 17496 21180 17524
rect 21174 17484 21180 17496
rect 21232 17484 21238 17536
rect 22005 17527 22063 17533
rect 22005 17493 22017 17527
rect 22051 17524 22063 17527
rect 22738 17524 22744 17536
rect 22051 17496 22744 17524
rect 22051 17493 22063 17496
rect 22005 17487 22063 17493
rect 22738 17484 22744 17496
rect 22796 17484 22802 17536
rect 23216 17533 23244 17632
rect 23382 17620 23388 17672
rect 23440 17660 23446 17672
rect 23860 17660 23888 17691
rect 25130 17688 25136 17700
rect 25188 17688 25194 17740
rect 25222 17688 25228 17740
rect 25280 17728 25286 17740
rect 25516 17737 25544 17768
rect 35161 17765 35173 17799
rect 35207 17765 35219 17799
rect 35161 17759 35219 17765
rect 25317 17731 25375 17737
rect 25317 17728 25329 17731
rect 25280 17700 25329 17728
rect 25280 17688 25286 17700
rect 25317 17697 25329 17700
rect 25363 17697 25375 17731
rect 25317 17691 25375 17697
rect 25501 17731 25559 17737
rect 25501 17697 25513 17731
rect 25547 17697 25559 17731
rect 26694 17728 26700 17740
rect 26655 17700 26700 17728
rect 25501 17691 25559 17697
rect 26694 17688 26700 17700
rect 26752 17688 26758 17740
rect 30009 17731 30067 17737
rect 30009 17697 30021 17731
rect 30055 17728 30067 17731
rect 30374 17728 30380 17740
rect 30055 17700 30380 17728
rect 30055 17697 30067 17700
rect 30009 17691 30067 17697
rect 30374 17688 30380 17700
rect 30432 17688 30438 17740
rect 31202 17728 31208 17740
rect 31163 17700 31208 17728
rect 31202 17688 31208 17700
rect 31260 17688 31266 17740
rect 32674 17688 32680 17740
rect 32732 17728 32738 17740
rect 33505 17731 33563 17737
rect 33505 17728 33517 17731
rect 32732 17700 33517 17728
rect 32732 17688 32738 17700
rect 33505 17697 33517 17700
rect 33551 17728 33563 17731
rect 34790 17728 34796 17740
rect 33551 17700 34796 17728
rect 33551 17697 33563 17700
rect 33505 17691 33563 17697
rect 34790 17688 34796 17700
rect 34848 17728 34854 17740
rect 34848 17700 34928 17728
rect 34848 17688 34854 17700
rect 23440 17632 23888 17660
rect 24581 17663 24639 17669
rect 23440 17620 23446 17632
rect 24581 17629 24593 17663
rect 24627 17660 24639 17663
rect 25406 17660 25412 17672
rect 24627 17632 25412 17660
rect 24627 17629 24639 17632
rect 24581 17623 24639 17629
rect 25406 17620 25412 17632
rect 25464 17620 25470 17672
rect 26418 17660 26424 17672
rect 26379 17632 26424 17660
rect 26418 17620 26424 17632
rect 26476 17620 26482 17672
rect 27798 17620 27804 17672
rect 27856 17620 27862 17672
rect 28813 17663 28871 17669
rect 28813 17629 28825 17663
rect 28859 17660 28871 17663
rect 28902 17660 28908 17672
rect 28859 17632 28908 17660
rect 28859 17629 28871 17632
rect 28813 17623 28871 17629
rect 28902 17620 28908 17632
rect 28960 17620 28966 17672
rect 28997 17663 29055 17669
rect 28997 17629 29009 17663
rect 29043 17660 29055 17663
rect 29178 17660 29184 17672
rect 29043 17632 29184 17660
rect 29043 17629 29055 17632
rect 28997 17623 29055 17629
rect 29178 17620 29184 17632
rect 29236 17620 29242 17672
rect 29914 17660 29920 17672
rect 29875 17632 29920 17660
rect 29914 17620 29920 17632
rect 29972 17620 29978 17672
rect 32950 17660 32956 17672
rect 32911 17632 32956 17660
rect 32950 17620 32956 17632
rect 33008 17620 33014 17672
rect 33597 17663 33655 17669
rect 33597 17629 33609 17663
rect 33643 17660 33655 17663
rect 34054 17660 34060 17672
rect 33643 17632 34060 17660
rect 33643 17629 33655 17632
rect 33597 17623 33655 17629
rect 34054 17620 34060 17632
rect 34112 17620 34118 17672
rect 34900 17669 34928 17700
rect 34885 17663 34943 17669
rect 34885 17629 34897 17663
rect 34931 17629 34943 17663
rect 35176 17660 35204 17759
rect 35621 17663 35679 17669
rect 35621 17660 35633 17663
rect 35176 17632 35633 17660
rect 34885 17623 34943 17629
rect 35621 17629 35633 17632
rect 35667 17629 35679 17663
rect 35621 17623 35679 17629
rect 35805 17663 35863 17669
rect 35805 17629 35817 17663
rect 35851 17629 35863 17663
rect 35805 17623 35863 17629
rect 23569 17595 23627 17601
rect 23569 17561 23581 17595
rect 23615 17592 23627 17595
rect 24854 17592 24860 17604
rect 23615 17564 24860 17592
rect 23615 17561 23627 17564
rect 23569 17555 23627 17561
rect 24854 17552 24860 17564
rect 24912 17552 24918 17604
rect 25314 17552 25320 17604
rect 25372 17592 25378 17604
rect 25593 17595 25651 17601
rect 25593 17592 25605 17595
rect 25372 17564 25605 17592
rect 25372 17552 25378 17564
rect 25593 17561 25605 17564
rect 25639 17561 25651 17595
rect 34072 17592 34100 17620
rect 34977 17595 35035 17601
rect 34977 17592 34989 17595
rect 34072 17564 34989 17592
rect 25593 17555 25651 17561
rect 34977 17561 34989 17564
rect 35023 17561 35035 17595
rect 34977 17555 35035 17561
rect 23201 17527 23259 17533
rect 23201 17493 23213 17527
rect 23247 17493 23259 17527
rect 24762 17524 24768 17536
rect 24723 17496 24768 17524
rect 23201 17487 23259 17493
rect 24762 17484 24768 17496
rect 24820 17484 24826 17536
rect 25608 17524 25636 17555
rect 35066 17552 35072 17604
rect 35124 17592 35130 17604
rect 35161 17595 35219 17601
rect 35161 17592 35173 17595
rect 35124 17564 35173 17592
rect 35124 17552 35130 17564
rect 35161 17561 35173 17564
rect 35207 17561 35219 17595
rect 35161 17555 35219 17561
rect 35342 17552 35348 17604
rect 35400 17592 35406 17604
rect 35820 17592 35848 17623
rect 35400 17564 35848 17592
rect 35400 17552 35406 17564
rect 28166 17524 28172 17536
rect 25608 17496 28172 17524
rect 28166 17484 28172 17496
rect 28224 17484 28230 17536
rect 30282 17524 30288 17536
rect 30243 17496 30288 17524
rect 30282 17484 30288 17496
rect 30340 17484 30346 17536
rect 35250 17484 35256 17536
rect 35308 17524 35314 17536
rect 35713 17527 35771 17533
rect 35713 17524 35725 17527
rect 35308 17496 35725 17524
rect 35308 17484 35314 17496
rect 35713 17493 35725 17496
rect 35759 17493 35771 17527
rect 35713 17487 35771 17493
rect 1104 17434 37628 17456
rect 1104 17382 4874 17434
rect 4926 17382 4938 17434
rect 4990 17382 5002 17434
rect 5054 17382 5066 17434
rect 5118 17382 5130 17434
rect 5182 17382 35594 17434
rect 35646 17382 35658 17434
rect 35710 17382 35722 17434
rect 35774 17382 35786 17434
rect 35838 17382 35850 17434
rect 35902 17382 37628 17434
rect 1104 17360 37628 17382
rect 8202 17320 8208 17332
rect 1780 17292 8208 17320
rect 1780 17193 1808 17292
rect 8202 17280 8208 17292
rect 8260 17280 8266 17332
rect 8297 17323 8355 17329
rect 8297 17289 8309 17323
rect 8343 17289 8355 17323
rect 8754 17320 8760 17332
rect 8715 17292 8760 17320
rect 8297 17283 8355 17289
rect 5905 17255 5963 17261
rect 5905 17221 5917 17255
rect 5951 17252 5963 17255
rect 8312 17252 8340 17283
rect 8754 17280 8760 17292
rect 8812 17280 8818 17332
rect 9125 17323 9183 17329
rect 9125 17289 9137 17323
rect 9171 17320 9183 17323
rect 9674 17320 9680 17332
rect 9171 17292 9680 17320
rect 9171 17289 9183 17292
rect 9125 17283 9183 17289
rect 9674 17280 9680 17292
rect 9732 17320 9738 17332
rect 10413 17323 10471 17329
rect 10413 17320 10425 17323
rect 9732 17292 10425 17320
rect 9732 17280 9738 17292
rect 10413 17289 10425 17292
rect 10459 17289 10471 17323
rect 10413 17283 10471 17289
rect 10502 17280 10508 17332
rect 10560 17320 10566 17332
rect 11701 17323 11759 17329
rect 11701 17320 11713 17323
rect 10560 17292 11713 17320
rect 10560 17280 10566 17292
rect 11701 17289 11713 17292
rect 11747 17289 11759 17323
rect 12158 17320 12164 17332
rect 12119 17292 12164 17320
rect 11701 17283 11759 17289
rect 12158 17280 12164 17292
rect 12216 17280 12222 17332
rect 13630 17280 13636 17332
rect 13688 17320 13694 17332
rect 17221 17323 17279 17329
rect 13688 17292 16712 17320
rect 13688 17280 13694 17292
rect 10321 17255 10379 17261
rect 10321 17252 10333 17255
rect 5951 17224 7314 17252
rect 8312 17224 10333 17252
rect 5951 17221 5963 17224
rect 5905 17215 5963 17221
rect 1765 17187 1823 17193
rect 1765 17153 1777 17187
rect 1811 17153 1823 17187
rect 5810 17184 5816 17196
rect 5723 17156 5816 17184
rect 1765 17147 1823 17153
rect 5810 17144 5816 17156
rect 5868 17184 5874 17196
rect 6086 17184 6092 17196
rect 5868 17156 6092 17184
rect 5868 17144 5874 17156
rect 6086 17144 6092 17156
rect 6144 17144 6150 17196
rect 6546 17116 6552 17128
rect 6507 17088 6552 17116
rect 6546 17076 6552 17088
rect 6604 17076 6610 17128
rect 6822 17116 6828 17128
rect 6783 17088 6828 17116
rect 6822 17076 6828 17088
rect 6880 17076 6886 17128
rect 1578 16980 1584 16992
rect 1539 16952 1584 16980
rect 1578 16940 1584 16952
rect 1636 16940 1642 16992
rect 6822 16940 6828 16992
rect 6880 16980 6886 16992
rect 8312 16980 8340 17224
rect 10321 17221 10333 17224
rect 10367 17221 10379 17255
rect 10321 17215 10379 17221
rect 15562 17212 15568 17264
rect 15620 17212 15626 17264
rect 12069 17187 12127 17193
rect 12069 17153 12081 17187
rect 12115 17184 12127 17187
rect 12434 17184 12440 17196
rect 12115 17156 12440 17184
rect 12115 17153 12127 17156
rect 12069 17147 12127 17153
rect 12434 17144 12440 17156
rect 12492 17184 12498 17196
rect 13173 17187 13231 17193
rect 13173 17184 13185 17187
rect 12492 17156 13185 17184
rect 12492 17144 12498 17156
rect 13173 17153 13185 17156
rect 13219 17153 13231 17187
rect 13173 17147 13231 17153
rect 13265 17187 13323 17193
rect 13265 17153 13277 17187
rect 13311 17184 13323 17187
rect 14090 17184 14096 17196
rect 13311 17156 14096 17184
rect 13311 17153 13323 17156
rect 13265 17147 13323 17153
rect 14090 17144 14096 17156
rect 14148 17144 14154 17196
rect 9214 17116 9220 17128
rect 9175 17088 9220 17116
rect 9214 17076 9220 17088
rect 9272 17076 9278 17128
rect 9309 17119 9367 17125
rect 9309 17085 9321 17119
rect 9355 17085 9367 17119
rect 10594 17116 10600 17128
rect 10555 17088 10600 17116
rect 9309 17079 9367 17085
rect 9030 17008 9036 17060
rect 9088 17048 9094 17060
rect 9324 17048 9352 17079
rect 10594 17076 10600 17088
rect 10652 17076 10658 17128
rect 12345 17119 12403 17125
rect 12345 17085 12357 17119
rect 12391 17116 12403 17119
rect 12894 17116 12900 17128
rect 12391 17088 12900 17116
rect 12391 17085 12403 17088
rect 12345 17079 12403 17085
rect 12894 17076 12900 17088
rect 12952 17076 12958 17128
rect 13081 17119 13139 17125
rect 13081 17085 13093 17119
rect 13127 17116 13139 17119
rect 13354 17116 13360 17128
rect 13127 17088 13360 17116
rect 13127 17085 13139 17088
rect 13081 17079 13139 17085
rect 13354 17076 13360 17088
rect 13412 17076 13418 17128
rect 14553 17119 14611 17125
rect 14553 17085 14565 17119
rect 14599 17085 14611 17119
rect 14826 17116 14832 17128
rect 14787 17088 14832 17116
rect 14553 17079 14611 17085
rect 9088 17020 9352 17048
rect 9088 17008 9094 17020
rect 13262 17008 13268 17060
rect 13320 17048 13326 17060
rect 14568 17048 14596 17079
rect 14826 17076 14832 17088
rect 14884 17076 14890 17128
rect 15286 17076 15292 17128
rect 15344 17116 15350 17128
rect 16301 17119 16359 17125
rect 16301 17116 16313 17119
rect 15344 17088 16313 17116
rect 15344 17076 15350 17088
rect 16301 17085 16313 17088
rect 16347 17116 16359 17119
rect 16482 17116 16488 17128
rect 16347 17088 16488 17116
rect 16347 17085 16359 17088
rect 16301 17079 16359 17085
rect 16482 17076 16488 17088
rect 16540 17076 16546 17128
rect 16684 17116 16712 17292
rect 17221 17289 17233 17323
rect 17267 17320 17279 17323
rect 17586 17320 17592 17332
rect 17267 17292 17592 17320
rect 17267 17289 17279 17292
rect 17221 17283 17279 17289
rect 17586 17280 17592 17292
rect 17644 17280 17650 17332
rect 18874 17320 18880 17332
rect 18835 17292 18880 17320
rect 18874 17280 18880 17292
rect 18932 17280 18938 17332
rect 19705 17323 19763 17329
rect 19705 17289 19717 17323
rect 19751 17320 19763 17323
rect 21082 17320 21088 17332
rect 19751 17292 21088 17320
rect 19751 17289 19763 17292
rect 19705 17283 19763 17289
rect 21082 17280 21088 17292
rect 21140 17280 21146 17332
rect 23658 17280 23664 17332
rect 23716 17320 23722 17332
rect 24581 17323 24639 17329
rect 24581 17320 24593 17323
rect 23716 17292 24593 17320
rect 23716 17280 23722 17292
rect 24581 17289 24593 17292
rect 24627 17289 24639 17323
rect 25406 17320 25412 17332
rect 25367 17292 25412 17320
rect 24581 17283 24639 17289
rect 25406 17280 25412 17292
rect 25464 17280 25470 17332
rect 28261 17323 28319 17329
rect 28261 17289 28273 17323
rect 28307 17320 28319 17323
rect 28534 17320 28540 17332
rect 28307 17292 28540 17320
rect 28307 17289 28319 17292
rect 28261 17283 28319 17289
rect 28534 17280 28540 17292
rect 28592 17280 28598 17332
rect 29457 17323 29515 17329
rect 29457 17320 29469 17323
rect 28920 17292 29469 17320
rect 17313 17255 17371 17261
rect 17313 17221 17325 17255
rect 17359 17252 17371 17255
rect 17494 17252 17500 17264
rect 17359 17224 17500 17252
rect 17359 17221 17371 17224
rect 17313 17215 17371 17221
rect 17494 17212 17500 17224
rect 17552 17212 17558 17264
rect 20438 17212 20444 17264
rect 20496 17212 20502 17264
rect 21174 17252 21180 17264
rect 21135 17224 21180 17252
rect 21174 17212 21180 17224
rect 21232 17212 21238 17264
rect 22738 17212 22744 17264
rect 22796 17212 22802 17264
rect 28920 17261 28948 17292
rect 29457 17289 29469 17292
rect 29503 17320 29515 17323
rect 29914 17320 29920 17332
rect 29503 17292 29920 17320
rect 29503 17289 29515 17292
rect 29457 17283 29515 17289
rect 29914 17280 29920 17292
rect 29972 17280 29978 17332
rect 30374 17320 30380 17332
rect 30116 17292 30380 17320
rect 28813 17255 28871 17261
rect 28813 17252 28825 17255
rect 27264 17224 28825 17252
rect 27264 17196 27292 17224
rect 28813 17221 28825 17224
rect 28859 17221 28871 17255
rect 28813 17215 28871 17221
rect 28905 17255 28963 17261
rect 28905 17221 28917 17255
rect 28951 17221 28963 17255
rect 30116 17252 30144 17292
rect 30374 17280 30380 17292
rect 30432 17320 30438 17332
rect 31202 17320 31208 17332
rect 30432 17292 31208 17320
rect 30432 17280 30438 17292
rect 31202 17280 31208 17292
rect 31260 17320 31266 17332
rect 34330 17320 34336 17332
rect 31260 17292 34336 17320
rect 31260 17280 31266 17292
rect 30282 17252 30288 17264
rect 28905 17215 28963 17221
rect 30024 17224 30144 17252
rect 30243 17224 30288 17252
rect 24673 17187 24731 17193
rect 24673 17153 24685 17187
rect 24719 17184 24731 17187
rect 25777 17187 25835 17193
rect 25777 17184 25789 17187
rect 24719 17156 25789 17184
rect 24719 17153 24731 17156
rect 24673 17147 24731 17153
rect 25777 17153 25789 17156
rect 25823 17184 25835 17187
rect 27246 17184 27252 17196
rect 25823 17156 27252 17184
rect 25823 17153 25835 17156
rect 25777 17147 25835 17153
rect 27246 17144 27252 17156
rect 27304 17144 27310 17196
rect 27341 17187 27399 17193
rect 27341 17153 27353 17187
rect 27387 17153 27399 17187
rect 27341 17147 27399 17153
rect 28537 17187 28595 17193
rect 28537 17153 28549 17187
rect 28583 17184 28595 17187
rect 28994 17184 29000 17196
rect 28583 17156 29000 17184
rect 28583 17153 28595 17156
rect 28537 17147 28595 17153
rect 17405 17119 17463 17125
rect 17405 17116 17417 17119
rect 16684 17088 17417 17116
rect 17405 17085 17417 17088
rect 17451 17116 17463 17119
rect 18601 17119 18659 17125
rect 18601 17116 18613 17119
rect 17451 17088 18613 17116
rect 17451 17085 17463 17088
rect 17405 17079 17463 17085
rect 18601 17085 18613 17088
rect 18647 17116 18659 17119
rect 18690 17116 18696 17128
rect 18647 17088 18696 17116
rect 18647 17085 18659 17088
rect 18601 17079 18659 17085
rect 18690 17076 18696 17088
rect 18748 17076 18754 17128
rect 18785 17119 18843 17125
rect 18785 17085 18797 17119
rect 18831 17116 18843 17119
rect 20714 17116 20720 17128
rect 18831 17088 20720 17116
rect 18831 17085 18843 17088
rect 18785 17079 18843 17085
rect 20714 17076 20720 17088
rect 20772 17076 20778 17128
rect 21453 17119 21511 17125
rect 21453 17085 21465 17119
rect 21499 17116 21511 17119
rect 21634 17116 21640 17128
rect 21499 17088 21640 17116
rect 21499 17085 21511 17088
rect 21453 17079 21511 17085
rect 21634 17076 21640 17088
rect 21692 17116 21698 17128
rect 22002 17116 22008 17128
rect 21692 17088 22008 17116
rect 21692 17076 21698 17088
rect 22002 17076 22008 17088
rect 22060 17076 22066 17128
rect 22278 17116 22284 17128
rect 22239 17088 22284 17116
rect 22278 17076 22284 17088
rect 22336 17076 22342 17128
rect 24857 17119 24915 17125
rect 24857 17085 24869 17119
rect 24903 17116 24915 17119
rect 24946 17116 24952 17128
rect 24903 17088 24952 17116
rect 24903 17085 24915 17088
rect 24857 17079 24915 17085
rect 24946 17076 24952 17088
rect 25004 17116 25010 17128
rect 25498 17116 25504 17128
rect 25004 17088 25504 17116
rect 25004 17076 25010 17088
rect 25498 17076 25504 17088
rect 25556 17076 25562 17128
rect 25869 17119 25927 17125
rect 25869 17085 25881 17119
rect 25915 17085 25927 17119
rect 25869 17079 25927 17085
rect 25961 17119 26019 17125
rect 25961 17085 25973 17119
rect 26007 17085 26019 17119
rect 25961 17079 26019 17085
rect 16758 17048 16764 17060
rect 13320 17020 14596 17048
rect 13320 17008 13326 17020
rect 9950 16980 9956 16992
rect 6880 16952 8340 16980
rect 9911 16952 9956 16980
rect 6880 16940 6886 16952
rect 9950 16940 9956 16952
rect 10008 16940 10014 16992
rect 13630 16980 13636 16992
rect 13591 16952 13636 16980
rect 13630 16940 13636 16952
rect 13688 16940 13694 16992
rect 14568 16980 14596 17020
rect 16224 17020 16764 17048
rect 16224 16980 16252 17020
rect 16758 17008 16764 17020
rect 16816 17008 16822 17060
rect 23474 17008 23480 17060
rect 23532 17048 23538 17060
rect 23753 17051 23811 17057
rect 23753 17048 23765 17051
rect 23532 17020 23765 17048
rect 23532 17008 23538 17020
rect 23753 17017 23765 17020
rect 23799 17048 23811 17051
rect 24578 17048 24584 17060
rect 23799 17020 24584 17048
rect 23799 17017 23811 17020
rect 23753 17011 23811 17017
rect 24578 17008 24584 17020
rect 24636 17048 24642 17060
rect 25884 17048 25912 17079
rect 24636 17020 25912 17048
rect 24636 17008 24642 17020
rect 14568 16952 16252 16980
rect 16853 16983 16911 16989
rect 16853 16949 16865 16983
rect 16899 16980 16911 16983
rect 16942 16980 16948 16992
rect 16899 16952 16948 16980
rect 16899 16949 16911 16952
rect 16853 16943 16911 16949
rect 16942 16940 16948 16952
rect 17000 16940 17006 16992
rect 18874 16940 18880 16992
rect 18932 16980 18938 16992
rect 19245 16983 19303 16989
rect 19245 16980 19257 16983
rect 18932 16952 19257 16980
rect 18932 16940 18938 16952
rect 19245 16949 19257 16952
rect 19291 16949 19303 16983
rect 24210 16980 24216 16992
rect 24171 16952 24216 16980
rect 19245 16943 19303 16949
rect 24210 16940 24216 16952
rect 24268 16940 24274 16992
rect 25222 16940 25228 16992
rect 25280 16980 25286 16992
rect 25498 16980 25504 16992
rect 25280 16952 25504 16980
rect 25280 16940 25286 16952
rect 25498 16940 25504 16952
rect 25556 16980 25562 16992
rect 25976 16980 26004 17079
rect 27154 17076 27160 17128
rect 27212 17116 27218 17128
rect 27356 17116 27384 17147
rect 28994 17144 29000 17156
rect 29052 17144 29058 17196
rect 30024 17193 30052 17224
rect 30282 17212 30288 17224
rect 30340 17212 30346 17264
rect 31662 17252 31668 17264
rect 31510 17224 31668 17252
rect 31662 17212 31668 17224
rect 31720 17212 31726 17264
rect 32324 17193 32352 17292
rect 34330 17280 34336 17292
rect 34388 17280 34394 17332
rect 35066 17280 35072 17332
rect 35124 17320 35130 17332
rect 35434 17320 35440 17332
rect 35124 17292 35440 17320
rect 35124 17280 35130 17292
rect 35434 17280 35440 17292
rect 35492 17320 35498 17332
rect 36633 17323 36691 17329
rect 36633 17320 36645 17323
rect 35492 17292 36645 17320
rect 35492 17280 35498 17292
rect 36633 17289 36645 17292
rect 36679 17289 36691 17323
rect 36633 17283 36691 17289
rect 33226 17212 33232 17264
rect 33284 17212 33290 17264
rect 35161 17255 35219 17261
rect 35161 17221 35173 17255
rect 35207 17252 35219 17255
rect 35250 17252 35256 17264
rect 35207 17224 35256 17252
rect 35207 17221 35219 17224
rect 35161 17215 35219 17221
rect 35250 17212 35256 17224
rect 35308 17212 35314 17264
rect 35894 17212 35900 17264
rect 35952 17212 35958 17264
rect 29549 17187 29607 17193
rect 29549 17153 29561 17187
rect 29595 17153 29607 17187
rect 29549 17147 29607 17153
rect 30009 17187 30067 17193
rect 30009 17153 30021 17187
rect 30055 17153 30067 17187
rect 30009 17147 30067 17153
rect 32309 17187 32367 17193
rect 32309 17153 32321 17187
rect 32355 17153 32367 17187
rect 32309 17147 32367 17153
rect 27212 17088 27384 17116
rect 27212 17076 27218 17088
rect 28074 17076 28080 17128
rect 28132 17116 28138 17128
rect 28445 17119 28503 17125
rect 28445 17116 28457 17119
rect 28132 17088 28457 17116
rect 28132 17076 28138 17088
rect 28445 17085 28457 17088
rect 28491 17085 28503 17119
rect 28445 17079 28503 17085
rect 25556 16952 26004 16980
rect 25556 16940 25562 16952
rect 27062 16940 27068 16992
rect 27120 16980 27126 16992
rect 27249 16983 27307 16989
rect 27249 16980 27261 16983
rect 27120 16952 27261 16980
rect 27120 16940 27126 16952
rect 27249 16949 27261 16952
rect 27295 16949 27307 16983
rect 29564 16980 29592 17147
rect 34330 17144 34336 17196
rect 34388 17184 34394 17196
rect 34885 17187 34943 17193
rect 34885 17184 34897 17187
rect 34388 17156 34897 17184
rect 34388 17144 34394 17156
rect 34885 17153 34897 17156
rect 34931 17153 34943 17187
rect 34885 17147 34943 17153
rect 32585 17119 32643 17125
rect 32585 17085 32597 17119
rect 32631 17116 32643 17119
rect 33318 17116 33324 17128
rect 32631 17088 33324 17116
rect 32631 17085 32643 17088
rect 32585 17079 32643 17085
rect 33318 17076 33324 17088
rect 33376 17076 33382 17128
rect 34054 17116 34060 17128
rect 34015 17088 34060 17116
rect 34054 17076 34060 17088
rect 34112 17076 34118 17128
rect 31757 16983 31815 16989
rect 31757 16980 31769 16983
rect 29564 16952 31769 16980
rect 27249 16943 27307 16949
rect 31757 16949 31769 16952
rect 31803 16980 31815 16983
rect 31846 16980 31852 16992
rect 31803 16952 31852 16980
rect 31803 16949 31815 16952
rect 31757 16943 31815 16949
rect 31846 16940 31852 16952
rect 31904 16980 31910 16992
rect 32398 16980 32404 16992
rect 31904 16952 32404 16980
rect 31904 16940 31910 16952
rect 32398 16940 32404 16952
rect 32456 16940 32462 16992
rect 1104 16890 37628 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 37628 16890
rect 1104 16816 37628 16838
rect 7098 16736 7104 16788
rect 7156 16776 7162 16788
rect 9582 16776 9588 16788
rect 7156 16748 9588 16776
rect 7156 16736 7162 16748
rect 9582 16736 9588 16748
rect 9640 16776 9646 16788
rect 10686 16776 10692 16788
rect 9640 16748 10692 16776
rect 9640 16736 9646 16748
rect 10686 16736 10692 16748
rect 10744 16736 10750 16788
rect 13722 16736 13728 16788
rect 13780 16776 13786 16788
rect 14369 16779 14427 16785
rect 14369 16776 14381 16779
rect 13780 16748 14381 16776
rect 13780 16736 13786 16748
rect 14369 16745 14381 16748
rect 14415 16745 14427 16779
rect 18598 16776 18604 16788
rect 18559 16748 18604 16776
rect 14369 16739 14427 16745
rect 18598 16736 18604 16748
rect 18656 16736 18662 16788
rect 20714 16736 20720 16788
rect 20772 16776 20778 16788
rect 21177 16779 21235 16785
rect 21177 16776 21189 16779
rect 20772 16748 21189 16776
rect 20772 16736 20778 16748
rect 21177 16745 21189 16748
rect 21223 16745 21235 16779
rect 22278 16776 22284 16788
rect 22239 16748 22284 16776
rect 21177 16739 21235 16745
rect 22278 16736 22284 16748
rect 22336 16736 22342 16788
rect 24762 16736 24768 16788
rect 24820 16776 24826 16788
rect 25758 16779 25816 16785
rect 25758 16776 25770 16779
rect 24820 16748 25770 16776
rect 24820 16736 24826 16748
rect 25758 16745 25770 16748
rect 25804 16745 25816 16779
rect 27246 16776 27252 16788
rect 27207 16748 27252 16776
rect 25758 16739 25816 16745
rect 27246 16736 27252 16748
rect 27304 16776 27310 16788
rect 27614 16776 27620 16788
rect 27304 16748 27620 16776
rect 27304 16736 27310 16748
rect 27614 16736 27620 16748
rect 27672 16736 27678 16788
rect 29178 16736 29184 16788
rect 29236 16776 29242 16788
rect 29825 16779 29883 16785
rect 29825 16776 29837 16779
rect 29236 16748 29837 16776
rect 29236 16736 29242 16748
rect 29825 16745 29837 16748
rect 29871 16745 29883 16779
rect 30742 16776 30748 16788
rect 30703 16748 30748 16776
rect 29825 16739 29883 16745
rect 30742 16736 30748 16748
rect 30800 16736 30806 16788
rect 30926 16776 30932 16788
rect 30887 16748 30932 16776
rect 30926 16736 30932 16748
rect 30984 16736 30990 16788
rect 34790 16736 34796 16788
rect 34848 16776 34854 16788
rect 35069 16779 35127 16785
rect 35069 16776 35081 16779
rect 34848 16748 35081 16776
rect 34848 16736 34854 16748
rect 35069 16745 35081 16748
rect 35115 16745 35127 16779
rect 35069 16739 35127 16745
rect 35253 16779 35311 16785
rect 35253 16745 35265 16779
rect 35299 16776 35311 16779
rect 35342 16776 35348 16788
rect 35299 16748 35348 16776
rect 35299 16745 35311 16748
rect 35253 16739 35311 16745
rect 35342 16736 35348 16748
rect 35400 16736 35406 16788
rect 35894 16736 35900 16788
rect 35952 16776 35958 16788
rect 35989 16779 36047 16785
rect 35989 16776 36001 16779
rect 35952 16748 36001 16776
rect 35952 16736 35958 16748
rect 35989 16745 36001 16748
rect 36035 16745 36047 16779
rect 35989 16739 36047 16745
rect 6086 16668 6092 16720
rect 6144 16708 6150 16720
rect 14090 16708 14096 16720
rect 6144 16680 9168 16708
rect 6144 16668 6150 16680
rect 6822 16640 6828 16652
rect 6783 16612 6828 16640
rect 6822 16600 6828 16612
rect 6880 16600 6886 16652
rect 6917 16643 6975 16649
rect 6917 16609 6929 16643
rect 6963 16640 6975 16643
rect 7190 16640 7196 16652
rect 6963 16612 7196 16640
rect 6963 16609 6975 16612
rect 6917 16603 6975 16609
rect 7190 16600 7196 16612
rect 7248 16600 7254 16652
rect 8021 16643 8079 16649
rect 8021 16609 8033 16643
rect 8067 16609 8079 16643
rect 8202 16640 8208 16652
rect 8163 16612 8208 16640
rect 8021 16603 8079 16609
rect 6733 16575 6791 16581
rect 6733 16541 6745 16575
rect 6779 16572 6791 16575
rect 7006 16572 7012 16584
rect 6779 16544 7012 16572
rect 6779 16541 6791 16544
rect 6733 16535 6791 16541
rect 7006 16532 7012 16544
rect 7064 16572 7070 16584
rect 8036 16572 8064 16603
rect 8202 16600 8208 16612
rect 8260 16600 8266 16652
rect 9140 16649 9168 16680
rect 12728 16680 14096 16708
rect 12728 16649 12756 16680
rect 14090 16668 14096 16680
rect 14148 16668 14154 16720
rect 23382 16668 23388 16720
rect 23440 16708 23446 16720
rect 24946 16708 24952 16720
rect 23440 16680 23612 16708
rect 24907 16680 24952 16708
rect 23440 16668 23446 16680
rect 9125 16643 9183 16649
rect 9125 16609 9137 16643
rect 9171 16609 9183 16643
rect 9125 16603 9183 16609
rect 12713 16643 12771 16649
rect 12713 16609 12725 16643
rect 12759 16609 12771 16643
rect 12713 16603 12771 16609
rect 12894 16600 12900 16652
rect 12952 16640 12958 16652
rect 13354 16640 13360 16652
rect 12952 16612 13360 16640
rect 12952 16600 12958 16612
rect 13354 16600 13360 16612
rect 13412 16600 13418 16652
rect 14274 16600 14280 16652
rect 14332 16640 14338 16652
rect 14332 16612 16160 16640
rect 14332 16600 14338 16612
rect 7064 16544 8064 16572
rect 7064 16532 7070 16544
rect 10778 16532 10784 16584
rect 10836 16572 10842 16584
rect 11609 16575 11667 16581
rect 11609 16572 11621 16575
rect 10836 16544 11621 16572
rect 10836 16532 10842 16544
rect 11609 16541 11621 16544
rect 11655 16572 11667 16575
rect 13630 16572 13636 16584
rect 11655 16544 13492 16572
rect 13591 16544 13636 16572
rect 11655 16541 11667 16544
rect 11609 16535 11667 16541
rect 6638 16464 6644 16516
rect 6696 16504 6702 16516
rect 9398 16504 9404 16516
rect 6696 16476 7604 16504
rect 9359 16476 9404 16504
rect 6696 16464 6702 16476
rect 6362 16436 6368 16448
rect 6323 16408 6368 16436
rect 6362 16396 6368 16408
rect 6420 16396 6426 16448
rect 7576 16445 7604 16476
rect 9398 16464 9404 16476
rect 9456 16464 9462 16516
rect 10134 16464 10140 16516
rect 10192 16464 10198 16516
rect 12621 16507 12679 16513
rect 12621 16504 12633 16507
rect 10888 16476 12633 16504
rect 7561 16439 7619 16445
rect 7561 16405 7573 16439
rect 7607 16405 7619 16439
rect 7926 16436 7932 16448
rect 7887 16408 7932 16436
rect 7561 16399 7619 16405
rect 7926 16396 7932 16408
rect 7984 16396 7990 16448
rect 9214 16396 9220 16448
rect 9272 16436 9278 16448
rect 10888 16445 10916 16476
rect 12621 16473 12633 16476
rect 12667 16473 12679 16507
rect 13464 16504 13492 16544
rect 13630 16532 13636 16544
rect 13688 16532 13694 16584
rect 14642 16572 14648 16584
rect 14603 16544 14648 16572
rect 14642 16532 14648 16544
rect 14700 16532 14706 16584
rect 15473 16575 15531 16581
rect 15473 16541 15485 16575
rect 15519 16572 15531 16575
rect 15654 16572 15660 16584
rect 15519 16544 15660 16572
rect 15519 16541 15531 16544
rect 15473 16535 15531 16541
rect 15654 16532 15660 16544
rect 15712 16532 15718 16584
rect 16132 16581 16160 16612
rect 16758 16600 16764 16652
rect 16816 16640 16822 16652
rect 16853 16643 16911 16649
rect 16853 16640 16865 16643
rect 16816 16612 16865 16640
rect 16816 16600 16822 16612
rect 16853 16609 16865 16612
rect 16899 16609 16911 16643
rect 16853 16603 16911 16609
rect 19429 16643 19487 16649
rect 19429 16609 19441 16643
rect 19475 16640 19487 16643
rect 21634 16640 21640 16652
rect 19475 16612 21640 16640
rect 19475 16609 19487 16612
rect 19429 16603 19487 16609
rect 21634 16600 21640 16612
rect 21692 16600 21698 16652
rect 23474 16640 23480 16652
rect 23435 16612 23480 16640
rect 23474 16600 23480 16612
rect 23532 16600 23538 16652
rect 23584 16649 23612 16680
rect 24946 16668 24952 16680
rect 25004 16668 25010 16720
rect 28718 16708 28724 16720
rect 27908 16680 28724 16708
rect 23569 16643 23627 16649
rect 23569 16609 23581 16643
rect 23615 16609 23627 16643
rect 23569 16603 23627 16609
rect 25501 16643 25559 16649
rect 25501 16609 25513 16643
rect 25547 16640 25559 16643
rect 26418 16640 26424 16652
rect 25547 16612 26424 16640
rect 25547 16609 25559 16612
rect 25501 16603 25559 16609
rect 26418 16600 26424 16612
rect 26476 16600 26482 16652
rect 27154 16600 27160 16652
rect 27212 16640 27218 16652
rect 27908 16640 27936 16680
rect 28718 16668 28724 16680
rect 28776 16668 28782 16720
rect 28994 16668 29000 16720
rect 29052 16708 29058 16720
rect 32585 16711 32643 16717
rect 32585 16708 32597 16711
rect 29052 16680 32597 16708
rect 29052 16668 29058 16680
rect 32585 16677 32597 16680
rect 32631 16677 32643 16711
rect 32585 16671 32643 16677
rect 33428 16680 35940 16708
rect 33428 16652 33456 16680
rect 27212 16612 27936 16640
rect 27212 16600 27218 16612
rect 16117 16575 16175 16581
rect 16117 16541 16129 16575
rect 16163 16541 16175 16575
rect 16117 16535 16175 16541
rect 22097 16575 22155 16581
rect 22097 16541 22109 16575
rect 22143 16572 22155 16575
rect 23385 16575 23443 16581
rect 22143 16544 23060 16572
rect 22143 16541 22155 16544
rect 22097 16535 22155 16541
rect 14458 16504 14464 16516
rect 13464 16476 14464 16504
rect 12621 16467 12679 16473
rect 14458 16464 14464 16476
rect 14516 16464 14522 16516
rect 16574 16504 16580 16516
rect 15672 16476 16580 16504
rect 10873 16439 10931 16445
rect 10873 16436 10885 16439
rect 9272 16408 10885 16436
rect 9272 16396 9278 16408
rect 10873 16405 10885 16408
rect 10919 16405 10931 16439
rect 10873 16399 10931 16405
rect 11701 16439 11759 16445
rect 11701 16405 11713 16439
rect 11747 16436 11759 16439
rect 11974 16436 11980 16448
rect 11747 16408 11980 16436
rect 11747 16405 11759 16408
rect 11701 16399 11759 16405
rect 11974 16396 11980 16408
rect 12032 16396 12038 16448
rect 12250 16436 12256 16448
rect 12211 16408 12256 16436
rect 12250 16396 12256 16408
rect 12308 16396 12314 16448
rect 13449 16439 13507 16445
rect 13449 16405 13461 16439
rect 13495 16436 13507 16439
rect 13538 16436 13544 16448
rect 13495 16408 13544 16436
rect 13495 16405 13507 16408
rect 13449 16399 13507 16405
rect 13538 16396 13544 16408
rect 13596 16396 13602 16448
rect 15672 16445 15700 16476
rect 16574 16464 16580 16476
rect 16632 16464 16638 16516
rect 17126 16504 17132 16516
rect 17087 16476 17132 16504
rect 17126 16464 17132 16476
rect 17184 16464 17190 16516
rect 18138 16464 18144 16516
rect 18196 16464 18202 16516
rect 19334 16464 19340 16516
rect 19392 16504 19398 16516
rect 19705 16507 19763 16513
rect 19705 16504 19717 16507
rect 19392 16476 19717 16504
rect 19392 16464 19398 16476
rect 19705 16473 19717 16476
rect 19751 16473 19763 16507
rect 19705 16467 19763 16473
rect 20162 16464 20168 16516
rect 20220 16464 20226 16516
rect 15657 16439 15715 16445
rect 15657 16405 15669 16439
rect 15703 16405 15715 16439
rect 15657 16399 15715 16405
rect 16209 16439 16267 16445
rect 16209 16405 16221 16439
rect 16255 16436 16267 16439
rect 18046 16436 18052 16448
rect 16255 16408 18052 16436
rect 16255 16405 16267 16408
rect 16209 16399 16267 16405
rect 18046 16396 18052 16408
rect 18104 16396 18110 16448
rect 23032 16445 23060 16544
rect 23385 16541 23397 16575
rect 23431 16572 23443 16575
rect 24210 16572 24216 16584
rect 23431 16544 24216 16572
rect 23431 16541 23443 16544
rect 23385 16535 23443 16541
rect 24210 16532 24216 16544
rect 24268 16532 24274 16584
rect 27798 16572 27804 16584
rect 27759 16544 27804 16572
rect 27798 16532 27804 16544
rect 27856 16532 27862 16584
rect 27908 16581 27936 16612
rect 28166 16600 28172 16652
rect 28224 16640 28230 16652
rect 33410 16640 33416 16652
rect 28224 16612 28488 16640
rect 28224 16600 28230 16612
rect 28460 16581 28488 16612
rect 31772 16612 33416 16640
rect 27893 16575 27951 16581
rect 27893 16541 27905 16575
rect 27939 16541 27951 16575
rect 27893 16535 27951 16541
rect 28445 16575 28503 16581
rect 28445 16541 28457 16575
rect 28491 16541 28503 16575
rect 29730 16572 29736 16584
rect 29691 16544 29736 16572
rect 28445 16535 28503 16541
rect 29730 16532 29736 16544
rect 29788 16532 29794 16584
rect 30006 16572 30012 16584
rect 29967 16544 30012 16572
rect 30006 16532 30012 16544
rect 30064 16532 30070 16584
rect 31662 16572 31668 16584
rect 31623 16544 31668 16572
rect 31662 16532 31668 16544
rect 31720 16532 31726 16584
rect 31772 16581 31800 16612
rect 31757 16575 31815 16581
rect 31757 16541 31769 16575
rect 31803 16541 31815 16575
rect 32674 16572 32680 16584
rect 32635 16544 32680 16572
rect 31757 16535 31815 16541
rect 32674 16532 32680 16544
rect 32732 16532 32738 16584
rect 33060 16572 33088 16612
rect 33410 16600 33416 16612
rect 33468 16600 33474 16652
rect 34054 16640 34060 16652
rect 33980 16612 34060 16640
rect 33137 16575 33195 16581
rect 33137 16572 33149 16575
rect 33060 16544 33149 16572
rect 33137 16541 33149 16544
rect 33183 16541 33195 16575
rect 33137 16535 33195 16541
rect 33226 16532 33232 16584
rect 33284 16572 33290 16584
rect 33980 16581 34008 16612
rect 34054 16600 34060 16612
rect 34112 16640 34118 16652
rect 34112 16612 34928 16640
rect 34112 16600 34118 16612
rect 33965 16575 34023 16581
rect 33284 16544 33329 16572
rect 33284 16532 33290 16544
rect 33965 16541 33977 16575
rect 34011 16541 34023 16575
rect 33965 16535 34023 16541
rect 23106 16464 23112 16516
rect 23164 16504 23170 16516
rect 24486 16504 24492 16516
rect 23164 16476 24492 16504
rect 23164 16464 23170 16476
rect 24486 16464 24492 16476
rect 24544 16504 24550 16516
rect 24673 16507 24731 16513
rect 24673 16504 24685 16507
rect 24544 16476 24685 16504
rect 24544 16464 24550 16476
rect 24673 16473 24685 16476
rect 24719 16473 24731 16507
rect 27062 16504 27068 16516
rect 27002 16476 27068 16504
rect 24673 16467 24731 16473
rect 27062 16464 27068 16476
rect 27120 16464 27126 16516
rect 28626 16464 28632 16516
rect 28684 16504 28690 16516
rect 31113 16507 31171 16513
rect 31113 16504 31125 16507
rect 28684 16476 31125 16504
rect 28684 16464 28690 16476
rect 31113 16473 31125 16476
rect 31159 16504 31171 16507
rect 31846 16504 31852 16516
rect 31159 16476 31852 16504
rect 31159 16473 31171 16476
rect 31113 16467 31171 16473
rect 31846 16464 31852 16476
rect 31904 16464 31910 16516
rect 34900 16513 34928 16612
rect 35912 16581 35940 16680
rect 35897 16575 35955 16581
rect 35897 16541 35909 16575
rect 35943 16572 35955 16575
rect 36170 16572 36176 16584
rect 35943 16544 36176 16572
rect 35943 16541 35955 16544
rect 35897 16535 35955 16541
rect 36170 16532 36176 16544
rect 36228 16532 36234 16584
rect 36906 16572 36912 16584
rect 36867 16544 36912 16572
rect 36906 16532 36912 16544
rect 36964 16532 36970 16584
rect 34885 16507 34943 16513
rect 34885 16473 34897 16507
rect 34931 16473 34943 16507
rect 34885 16467 34943 16473
rect 35101 16507 35159 16513
rect 35101 16473 35113 16507
rect 35147 16504 35159 16507
rect 35434 16504 35440 16516
rect 35147 16476 35440 16504
rect 35147 16473 35159 16476
rect 35101 16467 35159 16473
rect 35434 16464 35440 16476
rect 35492 16464 35498 16516
rect 23017 16439 23075 16445
rect 23017 16405 23029 16439
rect 23063 16405 23075 16439
rect 23017 16399 23075 16405
rect 28537 16439 28595 16445
rect 28537 16405 28549 16439
rect 28583 16436 28595 16439
rect 28718 16436 28724 16448
rect 28583 16408 28724 16436
rect 28583 16405 28595 16408
rect 28537 16399 28595 16405
rect 28718 16396 28724 16408
rect 28776 16396 28782 16448
rect 30098 16396 30104 16448
rect 30156 16436 30162 16448
rect 30285 16439 30343 16445
rect 30285 16436 30297 16439
rect 30156 16408 30297 16436
rect 30156 16396 30162 16408
rect 30285 16405 30297 16408
rect 30331 16405 30343 16439
rect 30285 16399 30343 16405
rect 30466 16396 30472 16448
rect 30524 16436 30530 16448
rect 30903 16439 30961 16445
rect 30903 16436 30915 16439
rect 30524 16408 30915 16436
rect 30524 16396 30530 16408
rect 30903 16405 30915 16408
rect 30949 16405 30961 16439
rect 30903 16399 30961 16405
rect 33318 16396 33324 16448
rect 33376 16436 33382 16448
rect 33873 16439 33931 16445
rect 33873 16436 33885 16439
rect 33376 16408 33885 16436
rect 33376 16396 33382 16408
rect 33873 16405 33885 16408
rect 33919 16405 33931 16439
rect 37090 16436 37096 16448
rect 37051 16408 37096 16436
rect 33873 16399 33931 16405
rect 37090 16396 37096 16408
rect 37148 16396 37154 16448
rect 1104 16346 37628 16368
rect 1104 16294 4874 16346
rect 4926 16294 4938 16346
rect 4990 16294 5002 16346
rect 5054 16294 5066 16346
rect 5118 16294 5130 16346
rect 5182 16294 35594 16346
rect 35646 16294 35658 16346
rect 35710 16294 35722 16346
rect 35774 16294 35786 16346
rect 35838 16294 35850 16346
rect 35902 16294 37628 16346
rect 1104 16272 37628 16294
rect 1946 16192 1952 16244
rect 2004 16232 2010 16244
rect 6914 16232 6920 16244
rect 2004 16204 6920 16232
rect 2004 16192 2010 16204
rect 6914 16192 6920 16204
rect 6972 16232 6978 16244
rect 8113 16235 8171 16241
rect 6972 16204 7065 16232
rect 6972 16192 6978 16204
rect 8113 16201 8125 16235
rect 8159 16232 8171 16235
rect 9398 16232 9404 16244
rect 8159 16204 9404 16232
rect 8159 16201 8171 16204
rect 8113 16195 8171 16201
rect 9398 16192 9404 16204
rect 9456 16192 9462 16244
rect 10134 16192 10140 16244
rect 10192 16232 10198 16244
rect 10229 16235 10287 16241
rect 10229 16232 10241 16235
rect 10192 16204 10241 16232
rect 10192 16192 10198 16204
rect 10229 16201 10241 16204
rect 10275 16201 10287 16235
rect 10229 16195 10287 16201
rect 11701 16235 11759 16241
rect 11701 16201 11713 16235
rect 11747 16201 11759 16235
rect 11701 16195 11759 16201
rect 12069 16235 12127 16241
rect 12069 16201 12081 16235
rect 12115 16232 12127 16235
rect 12250 16232 12256 16244
rect 12115 16204 12256 16232
rect 12115 16201 12127 16204
rect 12069 16195 12127 16201
rect 8941 16167 8999 16173
rect 8941 16133 8953 16167
rect 8987 16164 8999 16167
rect 9950 16164 9956 16176
rect 8987 16136 9956 16164
rect 8987 16133 8999 16136
rect 8941 16127 8999 16133
rect 9950 16124 9956 16136
rect 10008 16124 10014 16176
rect 7009 16099 7067 16105
rect 7009 16065 7021 16099
rect 7055 16096 7067 16099
rect 7834 16096 7840 16108
rect 7055 16068 7840 16096
rect 7055 16065 7067 16068
rect 7009 16059 7067 16065
rect 7834 16056 7840 16068
rect 7892 16056 7898 16108
rect 7929 16099 7987 16105
rect 7929 16065 7941 16099
rect 7975 16096 7987 16099
rect 9033 16099 9091 16105
rect 7975 16068 8616 16096
rect 7975 16065 7987 16068
rect 7929 16059 7987 16065
rect 7190 16028 7196 16040
rect 7103 16000 7196 16028
rect 7190 15988 7196 16000
rect 7248 16028 7254 16040
rect 7248 16000 8524 16028
rect 7248 15988 7254 16000
rect 5534 15852 5540 15904
rect 5592 15892 5598 15904
rect 6549 15895 6607 15901
rect 6549 15892 6561 15895
rect 5592 15864 6561 15892
rect 5592 15852 5598 15864
rect 6549 15861 6561 15864
rect 6595 15861 6607 15895
rect 8496 15892 8524 16000
rect 8588 15969 8616 16068
rect 9033 16065 9045 16099
rect 9079 16096 9091 16099
rect 9214 16096 9220 16108
rect 9079 16068 9220 16096
rect 9079 16065 9091 16068
rect 9033 16059 9091 16065
rect 9214 16056 9220 16068
rect 9272 16056 9278 16108
rect 10137 16099 10195 16105
rect 10137 16065 10149 16099
rect 10183 16096 10195 16099
rect 10778 16096 10784 16108
rect 10183 16068 10784 16096
rect 10183 16065 10195 16068
rect 10137 16059 10195 16065
rect 10778 16056 10784 16068
rect 10836 16056 10842 16108
rect 10965 16099 11023 16105
rect 10965 16065 10977 16099
rect 11011 16096 11023 16099
rect 11716 16096 11744 16195
rect 12250 16192 12256 16204
rect 12308 16192 12314 16244
rect 13814 16192 13820 16244
rect 13872 16232 13878 16244
rect 13872 16204 15516 16232
rect 13872 16192 13878 16204
rect 13538 16164 13544 16176
rect 13499 16136 13544 16164
rect 13538 16124 13544 16136
rect 13596 16124 13602 16176
rect 15102 16164 15108 16176
rect 14766 16136 15108 16164
rect 15102 16124 15108 16136
rect 15160 16124 15166 16176
rect 15488 16164 15516 16204
rect 15562 16192 15568 16244
rect 15620 16232 15626 16244
rect 15657 16235 15715 16241
rect 15657 16232 15669 16235
rect 15620 16204 15669 16232
rect 15620 16192 15626 16204
rect 15657 16201 15669 16204
rect 15703 16201 15715 16235
rect 17126 16232 17132 16244
rect 17087 16204 17132 16232
rect 15657 16195 15715 16201
rect 17126 16192 17132 16204
rect 17184 16192 17190 16244
rect 18049 16235 18107 16241
rect 18049 16201 18061 16235
rect 18095 16232 18107 16235
rect 18138 16232 18144 16244
rect 18095 16204 18144 16232
rect 18095 16201 18107 16204
rect 18049 16195 18107 16201
rect 18138 16192 18144 16204
rect 18196 16192 18202 16244
rect 19061 16235 19119 16241
rect 19061 16201 19073 16235
rect 19107 16232 19119 16235
rect 19334 16232 19340 16244
rect 19107 16204 19340 16232
rect 19107 16201 19119 16204
rect 19061 16195 19119 16201
rect 19334 16192 19340 16204
rect 19392 16192 19398 16244
rect 19705 16235 19763 16241
rect 19705 16201 19717 16235
rect 19751 16232 19763 16235
rect 20162 16232 20168 16244
rect 19751 16204 20168 16232
rect 19751 16201 19763 16204
rect 19705 16195 19763 16201
rect 20162 16192 20168 16204
rect 20220 16192 20226 16244
rect 20349 16235 20407 16241
rect 20349 16201 20361 16235
rect 20395 16232 20407 16235
rect 20438 16232 20444 16244
rect 20395 16204 20444 16232
rect 20395 16201 20407 16204
rect 20349 16195 20407 16201
rect 20438 16192 20444 16204
rect 20496 16192 20502 16244
rect 23385 16235 23443 16241
rect 23385 16201 23397 16235
rect 23431 16232 23443 16235
rect 24213 16235 24271 16241
rect 24213 16232 24225 16235
rect 23431 16204 24225 16232
rect 23431 16201 23443 16204
rect 23385 16195 23443 16201
rect 24213 16201 24225 16204
rect 24259 16201 24271 16235
rect 24578 16232 24584 16244
rect 24539 16204 24584 16232
rect 24213 16195 24271 16201
rect 24578 16192 24584 16204
rect 24636 16192 24642 16244
rect 28810 16232 28816 16244
rect 28736 16204 28816 16232
rect 18230 16164 18236 16176
rect 15488 16136 18236 16164
rect 11011 16068 11744 16096
rect 12161 16099 12219 16105
rect 11011 16065 11023 16068
rect 10965 16059 11023 16065
rect 12161 16065 12173 16099
rect 12207 16096 12219 16099
rect 12434 16096 12440 16108
rect 12207 16068 12440 16096
rect 12207 16065 12219 16068
rect 12161 16059 12219 16065
rect 12434 16056 12440 16068
rect 12492 16096 12498 16108
rect 12986 16096 12992 16108
rect 12492 16068 12992 16096
rect 12492 16056 12498 16068
rect 12986 16056 12992 16068
rect 13044 16056 13050 16108
rect 15488 16096 15516 16136
rect 15565 16099 15623 16105
rect 15565 16096 15577 16099
rect 15488 16068 15577 16096
rect 15565 16065 15577 16068
rect 15611 16065 15623 16099
rect 16942 16096 16948 16108
rect 16903 16068 16948 16096
rect 15565 16059 15623 16065
rect 16942 16056 16948 16068
rect 17000 16056 17006 16108
rect 18156 16105 18184 16136
rect 18230 16124 18236 16136
rect 18288 16164 18294 16176
rect 23474 16164 23480 16176
rect 18288 16136 19656 16164
rect 23387 16136 23480 16164
rect 18288 16124 18294 16136
rect 18141 16099 18199 16105
rect 18141 16065 18153 16099
rect 18187 16065 18199 16099
rect 18874 16096 18880 16108
rect 18835 16068 18880 16096
rect 18141 16059 18199 16065
rect 18874 16056 18880 16068
rect 18932 16056 18938 16108
rect 19628 16105 19656 16136
rect 23474 16124 23480 16136
rect 23532 16164 23538 16176
rect 25685 16167 25743 16173
rect 25685 16164 25697 16167
rect 23532 16136 25697 16164
rect 23532 16124 23538 16136
rect 25685 16133 25697 16136
rect 25731 16133 25743 16167
rect 28626 16164 28632 16176
rect 28587 16136 28632 16164
rect 25685 16127 25743 16133
rect 28626 16124 28632 16136
rect 28684 16124 28690 16176
rect 28736 16173 28764 16204
rect 28810 16192 28816 16204
rect 28868 16192 28874 16244
rect 30006 16232 30012 16244
rect 29967 16204 30012 16232
rect 30006 16192 30012 16204
rect 30064 16192 30070 16244
rect 28721 16167 28779 16173
rect 28721 16133 28733 16167
rect 28767 16133 28779 16167
rect 31389 16167 31447 16173
rect 31389 16164 31401 16167
rect 28721 16127 28779 16133
rect 29288 16136 29960 16164
rect 19613 16099 19671 16105
rect 19613 16065 19625 16099
rect 19659 16096 19671 16099
rect 20257 16099 20315 16105
rect 20257 16096 20269 16099
rect 19659 16068 20269 16096
rect 19659 16065 19671 16068
rect 19613 16059 19671 16065
rect 20257 16065 20269 16068
rect 20303 16065 20315 16099
rect 20257 16059 20315 16065
rect 22373 16099 22431 16105
rect 22373 16065 22385 16099
rect 22419 16096 22431 16099
rect 24673 16099 24731 16105
rect 22419 16068 23060 16096
rect 22419 16065 22431 16068
rect 22373 16059 22431 16065
rect 9122 16028 9128 16040
rect 9083 16000 9128 16028
rect 9122 15988 9128 16000
rect 9180 16028 9186 16040
rect 9582 16028 9588 16040
rect 9180 16000 9588 16028
rect 9180 15988 9186 16000
rect 9582 15988 9588 16000
rect 9640 16028 9646 16040
rect 12253 16031 12311 16037
rect 12253 16028 12265 16031
rect 9640 16000 12265 16028
rect 9640 15988 9646 16000
rect 12253 15997 12265 16000
rect 12299 16028 12311 16031
rect 13078 16028 13084 16040
rect 12299 16000 13084 16028
rect 12299 15997 12311 16000
rect 12253 15991 12311 15997
rect 13078 15988 13084 16000
rect 13136 15988 13142 16040
rect 13262 16028 13268 16040
rect 13223 16000 13268 16028
rect 13262 15988 13268 16000
rect 13320 15988 13326 16040
rect 14090 15988 14096 16040
rect 14148 16028 14154 16040
rect 15013 16031 15071 16037
rect 15013 16028 15025 16031
rect 14148 16000 15025 16028
rect 14148 15988 14154 16000
rect 15013 15997 15025 16000
rect 15059 16028 15071 16031
rect 17954 16028 17960 16040
rect 15059 16000 17960 16028
rect 15059 15997 15071 16000
rect 15013 15991 15071 15997
rect 17954 15988 17960 16000
rect 18012 15988 18018 16040
rect 8573 15963 8631 15969
rect 8573 15929 8585 15963
rect 8619 15929 8631 15963
rect 8573 15923 8631 15929
rect 15194 15920 15200 15972
rect 15252 15960 15258 15972
rect 23032 15969 23060 16068
rect 24673 16065 24685 16099
rect 24719 16096 24731 16099
rect 25590 16096 25596 16108
rect 24719 16068 25596 16096
rect 24719 16065 24731 16068
rect 24673 16059 24731 16065
rect 25590 16056 25596 16068
rect 25648 16096 25654 16108
rect 25777 16099 25835 16105
rect 25777 16096 25789 16099
rect 25648 16068 25789 16096
rect 25648 16056 25654 16068
rect 25777 16065 25789 16068
rect 25823 16065 25835 16099
rect 25777 16059 25835 16065
rect 27154 16056 27160 16108
rect 27212 16096 27218 16108
rect 27341 16099 27399 16105
rect 27341 16096 27353 16099
rect 27212 16068 27353 16096
rect 27212 16056 27218 16068
rect 27341 16065 27353 16068
rect 27387 16065 27399 16099
rect 27341 16059 27399 16065
rect 27706 16056 27712 16108
rect 27764 16096 27770 16108
rect 28353 16099 28411 16105
rect 28353 16096 28365 16099
rect 27764 16068 28365 16096
rect 27764 16056 27770 16068
rect 28353 16065 28365 16068
rect 28399 16065 28411 16099
rect 28353 16059 28411 16065
rect 28442 16056 28448 16108
rect 28500 16096 28506 16108
rect 28859 16099 28917 16105
rect 28859 16096 28871 16099
rect 28500 16068 28545 16096
rect 28644 16068 28871 16096
rect 28500 16056 28506 16068
rect 28644 16040 28672 16068
rect 28859 16065 28871 16068
rect 28905 16096 28917 16099
rect 29288 16096 29316 16136
rect 29454 16096 29460 16108
rect 28905 16068 29316 16096
rect 29415 16068 29460 16096
rect 28905 16065 28917 16068
rect 28859 16059 28917 16065
rect 29454 16056 29460 16068
rect 29512 16056 29518 16108
rect 29546 16056 29552 16108
rect 29604 16096 29610 16108
rect 29733 16099 29791 16105
rect 29604 16068 29649 16096
rect 29604 16056 29610 16068
rect 29733 16065 29745 16099
rect 29779 16065 29791 16099
rect 29733 16059 29791 16065
rect 29825 16099 29883 16105
rect 29825 16065 29837 16099
rect 29871 16065 29883 16099
rect 29825 16059 29883 16065
rect 23382 15988 23388 16040
rect 23440 16028 23446 16040
rect 23569 16031 23627 16037
rect 23569 16028 23581 16031
rect 23440 16000 23581 16028
rect 23440 15988 23446 16000
rect 23569 15997 23581 16000
rect 23615 15997 23627 16031
rect 24762 16028 24768 16040
rect 24723 16000 24768 16028
rect 23569 15991 23627 15997
rect 24762 15988 24768 16000
rect 24820 15988 24826 16040
rect 25498 16028 25504 16040
rect 25459 16000 25504 16028
rect 25498 15988 25504 16000
rect 25556 15988 25562 16040
rect 28626 15988 28632 16040
rect 28684 15988 28690 16040
rect 29748 16028 29776 16059
rect 28736 16000 29776 16028
rect 28736 15972 28764 16000
rect 23017 15963 23075 15969
rect 15252 15932 22968 15960
rect 15252 15920 15258 15932
rect 9030 15892 9036 15904
rect 8496 15864 9036 15892
rect 6549 15855 6607 15861
rect 9030 15852 9036 15864
rect 9088 15892 9094 15904
rect 9398 15892 9404 15904
rect 9088 15864 9404 15892
rect 9088 15852 9094 15864
rect 9398 15852 9404 15864
rect 9456 15852 9462 15904
rect 11146 15892 11152 15904
rect 11107 15864 11152 15892
rect 11146 15852 11152 15864
rect 11204 15852 11210 15904
rect 21910 15852 21916 15904
rect 21968 15892 21974 15904
rect 22189 15895 22247 15901
rect 22189 15892 22201 15895
rect 21968 15864 22201 15892
rect 21968 15852 21974 15864
rect 22189 15861 22201 15864
rect 22235 15861 22247 15895
rect 22940 15892 22968 15932
rect 23017 15929 23029 15963
rect 23063 15929 23075 15963
rect 23017 15923 23075 15929
rect 26145 15963 26203 15969
rect 26145 15929 26157 15963
rect 26191 15960 26203 15963
rect 28534 15960 28540 15972
rect 26191 15932 28540 15960
rect 26191 15929 26203 15932
rect 26145 15923 26203 15929
rect 28534 15920 28540 15932
rect 28592 15920 28598 15972
rect 28718 15920 28724 15972
rect 28776 15920 28782 15972
rect 29840 15960 29868 16059
rect 29932 16028 29960 16136
rect 30852 16136 31401 16164
rect 30466 16056 30472 16108
rect 30524 16096 30530 16108
rect 30852 16105 30880 16136
rect 31389 16133 31401 16136
rect 31435 16133 31447 16167
rect 31389 16127 31447 16133
rect 32585 16167 32643 16173
rect 32585 16133 32597 16167
rect 32631 16164 32643 16167
rect 32766 16164 32772 16176
rect 32631 16136 32772 16164
rect 32631 16133 32643 16136
rect 32585 16127 32643 16133
rect 32766 16124 32772 16136
rect 32824 16124 32830 16176
rect 35434 16164 35440 16176
rect 34072 16136 35440 16164
rect 30653 16099 30711 16105
rect 30653 16096 30665 16099
rect 30524 16068 30665 16096
rect 30524 16056 30530 16068
rect 30653 16065 30665 16068
rect 30699 16065 30711 16099
rect 30653 16059 30711 16065
rect 30837 16099 30895 16105
rect 30837 16065 30849 16099
rect 30883 16065 30895 16099
rect 30837 16059 30895 16065
rect 30926 16056 30932 16108
rect 30984 16096 30990 16108
rect 31297 16099 31355 16105
rect 31297 16096 31309 16099
rect 30984 16068 31309 16096
rect 30984 16056 30990 16068
rect 31297 16065 31309 16068
rect 31343 16065 31355 16099
rect 31478 16096 31484 16108
rect 31439 16068 31484 16096
rect 31297 16059 31355 16065
rect 31478 16056 31484 16068
rect 31536 16056 31542 16108
rect 32401 16099 32459 16105
rect 32401 16065 32413 16099
rect 32447 16096 32459 16099
rect 32490 16096 32496 16108
rect 32447 16068 32496 16096
rect 32447 16065 32459 16068
rect 32401 16059 32459 16065
rect 32490 16056 32496 16068
rect 32548 16056 32554 16108
rect 32674 16056 32680 16108
rect 32732 16096 32738 16108
rect 34072 16105 34100 16136
rect 35434 16124 35440 16136
rect 35492 16124 35498 16176
rect 34057 16099 34115 16105
rect 32732 16068 32777 16096
rect 32732 16056 32738 16068
rect 34057 16065 34069 16099
rect 34103 16065 34115 16099
rect 34057 16059 34115 16065
rect 34701 16099 34759 16105
rect 34701 16065 34713 16099
rect 34747 16096 34759 16099
rect 35342 16096 35348 16108
rect 34747 16068 35348 16096
rect 34747 16065 34759 16068
rect 34701 16059 34759 16065
rect 35342 16056 35348 16068
rect 35400 16056 35406 16108
rect 35529 16099 35587 16105
rect 35529 16065 35541 16099
rect 35575 16065 35587 16099
rect 36170 16096 36176 16108
rect 36131 16068 36176 16096
rect 35529 16059 35587 16065
rect 34514 16028 34520 16040
rect 29932 16000 31754 16028
rect 34475 16000 34520 16028
rect 30742 15960 30748 15972
rect 29840 15932 30748 15960
rect 30742 15920 30748 15932
rect 30800 15920 30806 15972
rect 31726 15960 31754 16000
rect 34514 15988 34520 16000
rect 34572 16028 34578 16040
rect 35544 16028 35572 16059
rect 36170 16056 36176 16068
rect 36228 16096 36234 16108
rect 36633 16099 36691 16105
rect 36633 16096 36645 16099
rect 36228 16068 36645 16096
rect 36228 16056 36234 16068
rect 36633 16065 36645 16068
rect 36679 16065 36691 16099
rect 36633 16059 36691 16065
rect 34572 16000 35572 16028
rect 34572 15988 34578 16000
rect 33965 15963 34023 15969
rect 33965 15960 33977 15963
rect 31726 15932 33977 15960
rect 33965 15929 33977 15932
rect 34011 15929 34023 15963
rect 33965 15923 34023 15929
rect 34606 15920 34612 15972
rect 34664 15960 34670 15972
rect 35345 15963 35403 15969
rect 35345 15960 35357 15963
rect 34664 15932 35357 15960
rect 34664 15920 34670 15932
rect 35345 15929 35357 15932
rect 35391 15929 35403 15963
rect 35345 15923 35403 15929
rect 23106 15892 23112 15904
rect 22940 15864 23112 15892
rect 22189 15855 22247 15861
rect 23106 15852 23112 15864
rect 23164 15852 23170 15904
rect 26602 15852 26608 15904
rect 26660 15892 26666 15904
rect 27249 15895 27307 15901
rect 27249 15892 27261 15895
rect 26660 15864 27261 15892
rect 26660 15852 26666 15864
rect 27249 15861 27261 15864
rect 27295 15861 27307 15895
rect 28994 15892 29000 15904
rect 28955 15864 29000 15892
rect 27249 15855 27307 15861
rect 28994 15852 29000 15864
rect 29052 15852 29058 15904
rect 30650 15852 30656 15904
rect 30708 15892 30714 15904
rect 30837 15895 30895 15901
rect 30837 15892 30849 15895
rect 30708 15864 30849 15892
rect 30708 15852 30714 15864
rect 30837 15861 30849 15864
rect 30883 15861 30895 15895
rect 32398 15892 32404 15904
rect 32359 15864 32404 15892
rect 30837 15855 30895 15861
rect 32398 15852 32404 15864
rect 32456 15852 32462 15904
rect 34790 15852 34796 15904
rect 34848 15892 34854 15904
rect 34885 15895 34943 15901
rect 34885 15892 34897 15895
rect 34848 15864 34897 15892
rect 34848 15852 34854 15864
rect 34885 15861 34897 15864
rect 34931 15861 34943 15895
rect 36078 15892 36084 15904
rect 36039 15864 36084 15892
rect 34885 15855 34943 15861
rect 36078 15852 36084 15864
rect 36136 15852 36142 15904
rect 36722 15892 36728 15904
rect 36683 15864 36728 15892
rect 36722 15852 36728 15864
rect 36780 15852 36786 15904
rect 1104 15802 37628 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 37628 15802
rect 1104 15728 37628 15750
rect 7926 15648 7932 15700
rect 7984 15688 7990 15700
rect 8021 15691 8079 15697
rect 8021 15688 8033 15691
rect 7984 15660 8033 15688
rect 7984 15648 7990 15660
rect 8021 15657 8033 15660
rect 8067 15657 8079 15691
rect 8021 15651 8079 15657
rect 11146 15648 11152 15700
rect 11204 15688 11210 15700
rect 11498 15691 11556 15697
rect 11498 15688 11510 15691
rect 11204 15660 11510 15688
rect 11204 15648 11210 15660
rect 11498 15657 11510 15660
rect 11544 15657 11556 15691
rect 12986 15688 12992 15700
rect 12947 15660 12992 15688
rect 11498 15651 11556 15657
rect 12986 15648 12992 15660
rect 13044 15648 13050 15700
rect 14826 15648 14832 15700
rect 14884 15688 14890 15700
rect 15197 15691 15255 15697
rect 15197 15688 15209 15691
rect 14884 15660 15209 15688
rect 14884 15648 14890 15660
rect 15197 15657 15209 15660
rect 15243 15657 15255 15691
rect 23385 15691 23443 15697
rect 15197 15651 15255 15657
rect 15948 15660 23336 15688
rect 8956 15592 11284 15620
rect 8956 15564 8984 15592
rect 6273 15555 6331 15561
rect 6273 15521 6285 15555
rect 6319 15552 6331 15555
rect 6546 15552 6552 15564
rect 6319 15524 6552 15552
rect 6319 15521 6331 15524
rect 6273 15515 6331 15521
rect 6546 15512 6552 15524
rect 6604 15552 6610 15564
rect 8294 15552 8300 15564
rect 6604 15524 8300 15552
rect 6604 15512 6610 15524
rect 8294 15512 8300 15524
rect 8352 15552 8358 15564
rect 8938 15552 8944 15564
rect 8352 15524 8944 15552
rect 8352 15512 8358 15524
rect 8938 15512 8944 15524
rect 8996 15512 9002 15564
rect 9398 15512 9404 15564
rect 9456 15552 9462 15564
rect 11256 15561 11284 15592
rect 13814 15580 13820 15632
rect 13872 15620 13878 15632
rect 14461 15623 14519 15629
rect 14461 15620 14473 15623
rect 13872 15592 14473 15620
rect 13872 15580 13878 15592
rect 14461 15589 14473 15592
rect 14507 15620 14519 15623
rect 15948 15620 15976 15660
rect 14507 15592 15976 15620
rect 23308 15620 23336 15660
rect 23385 15657 23397 15691
rect 23431 15688 23443 15691
rect 23474 15688 23480 15700
rect 23431 15660 23480 15688
rect 23431 15657 23443 15660
rect 23385 15651 23443 15657
rect 23474 15648 23480 15660
rect 23532 15648 23538 15700
rect 25041 15691 25099 15697
rect 25041 15657 25053 15691
rect 25087 15688 25099 15691
rect 25498 15688 25504 15700
rect 25087 15660 25504 15688
rect 25087 15657 25099 15660
rect 25041 15651 25099 15657
rect 25498 15648 25504 15660
rect 25556 15648 25562 15700
rect 27893 15691 27951 15697
rect 27893 15657 27905 15691
rect 27939 15688 27951 15691
rect 28442 15688 28448 15700
rect 27939 15660 28448 15688
rect 27939 15657 27951 15660
rect 27893 15651 27951 15657
rect 28442 15648 28448 15660
rect 28500 15648 28506 15700
rect 29181 15691 29239 15697
rect 29181 15657 29193 15691
rect 29227 15688 29239 15691
rect 29730 15688 29736 15700
rect 29227 15660 29736 15688
rect 29227 15657 29239 15660
rect 29181 15651 29239 15657
rect 29730 15648 29736 15660
rect 29788 15648 29794 15700
rect 29840 15660 31754 15688
rect 23842 15620 23848 15632
rect 23308 15592 23848 15620
rect 14507 15589 14519 15592
rect 14461 15583 14519 15589
rect 23842 15580 23848 15592
rect 23900 15580 23906 15632
rect 9677 15555 9735 15561
rect 9677 15552 9689 15555
rect 9456 15524 9689 15552
rect 9456 15512 9462 15524
rect 9677 15521 9689 15524
rect 9723 15521 9735 15555
rect 9677 15515 9735 15521
rect 11241 15555 11299 15561
rect 11241 15521 11253 15555
rect 11287 15552 11299 15555
rect 13262 15552 13268 15564
rect 11287 15524 13268 15552
rect 11287 15521 11299 15524
rect 11241 15515 11299 15521
rect 13262 15512 13268 15524
rect 13320 15512 13326 15564
rect 21910 15552 21916 15564
rect 21871 15524 21916 15552
rect 21910 15512 21916 15524
rect 21968 15512 21974 15564
rect 22646 15512 22652 15564
rect 22704 15552 22710 15564
rect 25866 15552 25872 15564
rect 22704 15524 25872 15552
rect 22704 15512 22710 15524
rect 5810 15484 5816 15496
rect 5771 15456 5816 15484
rect 5810 15444 5816 15456
rect 5868 15444 5874 15496
rect 8478 15444 8484 15496
rect 8536 15484 8542 15496
rect 9493 15487 9551 15493
rect 9493 15484 9505 15487
rect 8536 15456 9505 15484
rect 8536 15444 8542 15456
rect 9493 15453 9505 15456
rect 9539 15484 9551 15487
rect 9766 15484 9772 15496
rect 9539 15456 9772 15484
rect 9539 15453 9551 15456
rect 9493 15447 9551 15453
rect 9766 15444 9772 15456
rect 9824 15444 9830 15496
rect 9858 15444 9864 15496
rect 9916 15484 9922 15496
rect 10505 15487 10563 15493
rect 10505 15484 10517 15487
rect 9916 15456 10517 15484
rect 9916 15444 9922 15456
rect 10505 15453 10517 15456
rect 10551 15453 10563 15487
rect 10505 15447 10563 15453
rect 14645 15487 14703 15493
rect 14645 15453 14657 15487
rect 14691 15484 14703 15487
rect 15194 15484 15200 15496
rect 14691 15456 15200 15484
rect 14691 15453 14703 15456
rect 14645 15447 14703 15453
rect 6546 15416 6552 15428
rect 6507 15388 6552 15416
rect 6546 15376 6552 15388
rect 6604 15376 6610 15428
rect 6886 15388 7038 15416
rect 5721 15351 5779 15357
rect 5721 15317 5733 15351
rect 5767 15348 5779 15351
rect 6886 15348 6914 15388
rect 5767 15320 6914 15348
rect 5767 15317 5779 15320
rect 5721 15311 5779 15317
rect 8386 15308 8392 15360
rect 8444 15348 8450 15360
rect 9125 15351 9183 15357
rect 9125 15348 9137 15351
rect 8444 15320 9137 15348
rect 8444 15308 8450 15320
rect 9125 15317 9137 15320
rect 9171 15317 9183 15351
rect 9125 15311 9183 15317
rect 9585 15351 9643 15357
rect 9585 15317 9597 15351
rect 9631 15348 9643 15351
rect 10042 15348 10048 15360
rect 9631 15320 10048 15348
rect 9631 15317 9643 15320
rect 9585 15311 9643 15317
rect 10042 15308 10048 15320
rect 10100 15308 10106 15360
rect 10318 15308 10324 15360
rect 10376 15348 10382 15360
rect 10413 15351 10471 15357
rect 10413 15348 10425 15351
rect 10376 15320 10425 15348
rect 10376 15308 10382 15320
rect 10413 15317 10425 15320
rect 10459 15317 10471 15351
rect 10520 15348 10548 15447
rect 15194 15444 15200 15456
rect 15252 15444 15258 15496
rect 15378 15484 15384 15496
rect 15339 15456 15384 15484
rect 15378 15444 15384 15456
rect 15436 15444 15442 15496
rect 16301 15487 16359 15493
rect 16301 15453 16313 15487
rect 16347 15484 16359 15487
rect 17402 15484 17408 15496
rect 16347 15456 17408 15484
rect 16347 15453 16359 15456
rect 16301 15447 16359 15453
rect 17402 15444 17408 15456
rect 17460 15484 17466 15496
rect 18506 15484 18512 15496
rect 17460 15456 18512 15484
rect 17460 15444 17466 15456
rect 18506 15444 18512 15456
rect 18564 15444 18570 15496
rect 21634 15484 21640 15496
rect 21595 15456 21640 15484
rect 21634 15444 21640 15456
rect 21692 15444 21698 15496
rect 24780 15493 24808 15524
rect 25866 15512 25872 15524
rect 25924 15512 25930 15564
rect 28718 15552 28724 15564
rect 28679 15524 28724 15552
rect 28718 15512 28724 15524
rect 28776 15512 28782 15564
rect 28813 15555 28871 15561
rect 28813 15521 28825 15555
rect 28859 15552 28871 15555
rect 28902 15552 28908 15564
rect 28859 15524 28908 15552
rect 28859 15521 28871 15524
rect 28813 15515 28871 15521
rect 28902 15512 28908 15524
rect 28960 15552 28966 15564
rect 29840 15552 29868 15660
rect 31726 15620 31754 15660
rect 32490 15648 32496 15700
rect 32548 15688 32554 15700
rect 32585 15691 32643 15697
rect 32585 15688 32597 15691
rect 32548 15660 32597 15688
rect 32548 15648 32554 15660
rect 32585 15657 32597 15660
rect 32631 15657 32643 15691
rect 33318 15688 33324 15700
rect 32585 15651 32643 15657
rect 33060 15660 33324 15688
rect 33060 15620 33088 15660
rect 33318 15648 33324 15660
rect 33376 15648 33382 15700
rect 31726 15592 33088 15620
rect 30374 15552 30380 15564
rect 28960 15524 29868 15552
rect 30335 15524 30380 15552
rect 28960 15512 28966 15524
rect 30374 15512 30380 15524
rect 30432 15512 30438 15564
rect 30650 15552 30656 15564
rect 30611 15524 30656 15552
rect 30650 15512 30656 15524
rect 30708 15512 30714 15564
rect 34330 15552 34336 15564
rect 34291 15524 34336 15552
rect 34330 15512 34336 15524
rect 34388 15552 34394 15564
rect 35345 15555 35403 15561
rect 35345 15552 35357 15555
rect 34388 15524 35357 15552
rect 34388 15512 34394 15524
rect 35345 15521 35357 15524
rect 35391 15521 35403 15555
rect 35618 15552 35624 15564
rect 35579 15524 35624 15552
rect 35345 15515 35403 15521
rect 35618 15512 35624 15524
rect 35676 15512 35682 15564
rect 24765 15487 24823 15493
rect 24765 15453 24777 15487
rect 24811 15453 24823 15487
rect 24765 15447 24823 15453
rect 27338 15444 27344 15496
rect 27396 15484 27402 15496
rect 27396 15456 27441 15484
rect 27396 15444 27402 15456
rect 27614 15444 27620 15496
rect 27672 15484 27678 15496
rect 27801 15487 27859 15493
rect 27801 15484 27813 15487
rect 27672 15456 27813 15484
rect 27672 15444 27678 15456
rect 27801 15453 27813 15456
rect 27847 15453 27859 15487
rect 28442 15484 28448 15496
rect 28403 15456 28448 15484
rect 27801 15447 27859 15453
rect 28442 15444 28448 15456
rect 28500 15444 28506 15496
rect 28629 15487 28687 15493
rect 28629 15453 28641 15487
rect 28675 15453 28687 15487
rect 28629 15447 28687 15453
rect 28997 15487 29055 15493
rect 28997 15453 29009 15487
rect 29043 15484 29055 15487
rect 29454 15484 29460 15496
rect 29043 15456 29460 15484
rect 29043 15453 29055 15456
rect 28997 15447 29055 15453
rect 11974 15376 11980 15428
rect 12032 15376 12038 15428
rect 16025 15419 16083 15425
rect 12912 15388 14596 15416
rect 12912 15348 12940 15388
rect 10520 15320 12940 15348
rect 14568 15348 14596 15388
rect 16025 15385 16037 15419
rect 16071 15385 16083 15419
rect 16025 15379 16083 15385
rect 15378 15348 15384 15360
rect 14568 15320 15384 15348
rect 10413 15311 10471 15317
rect 15378 15308 15384 15320
rect 15436 15348 15442 15360
rect 16040 15348 16068 15379
rect 22646 15376 22652 15428
rect 22704 15376 22710 15428
rect 26602 15376 26608 15428
rect 26660 15376 26666 15428
rect 27062 15416 27068 15428
rect 27023 15388 27068 15416
rect 27062 15376 27068 15388
rect 27120 15376 27126 15428
rect 28644 15416 28672 15447
rect 29454 15444 29460 15456
rect 29512 15444 29518 15496
rect 29730 15484 29736 15496
rect 29691 15456 29736 15484
rect 29730 15444 29736 15456
rect 29788 15444 29794 15496
rect 29917 15487 29975 15493
rect 29917 15453 29929 15487
rect 29963 15484 29975 15487
rect 30282 15484 30288 15496
rect 29963 15456 30288 15484
rect 29963 15453 29975 15456
rect 29917 15447 29975 15453
rect 30282 15444 30288 15456
rect 30340 15444 30346 15496
rect 31754 15444 31760 15496
rect 31812 15444 31818 15496
rect 36722 15444 36728 15496
rect 36780 15444 36786 15496
rect 30742 15416 30748 15428
rect 28644 15388 30748 15416
rect 30742 15376 30748 15388
rect 30800 15376 30806 15428
rect 33042 15376 33048 15428
rect 33100 15376 33106 15428
rect 34054 15416 34060 15428
rect 34015 15388 34060 15416
rect 34054 15376 34060 15388
rect 34112 15376 34118 15428
rect 34164 15388 35756 15416
rect 25590 15348 25596 15360
rect 15436 15320 16068 15348
rect 25551 15320 25596 15348
rect 15436 15308 15442 15320
rect 25590 15308 25596 15320
rect 25648 15308 25654 15360
rect 29822 15348 29828 15360
rect 29783 15320 29828 15348
rect 29822 15308 29828 15320
rect 29880 15308 29886 15360
rect 30834 15308 30840 15360
rect 30892 15348 30898 15360
rect 31478 15348 31484 15360
rect 30892 15320 31484 15348
rect 30892 15308 30898 15320
rect 31478 15308 31484 15320
rect 31536 15348 31542 15360
rect 32125 15351 32183 15357
rect 32125 15348 32137 15351
rect 31536 15320 32137 15348
rect 31536 15308 31542 15320
rect 32125 15317 32137 15320
rect 32171 15317 32183 15351
rect 32125 15311 32183 15317
rect 32766 15308 32772 15360
rect 32824 15348 32830 15360
rect 34164 15348 34192 15388
rect 32824 15320 34192 15348
rect 35728 15348 35756 15388
rect 36262 15348 36268 15360
rect 35728 15320 36268 15348
rect 32824 15308 32830 15320
rect 36262 15308 36268 15320
rect 36320 15348 36326 15360
rect 37093 15351 37151 15357
rect 37093 15348 37105 15351
rect 36320 15320 37105 15348
rect 36320 15308 36326 15320
rect 37093 15317 37105 15320
rect 37139 15317 37151 15351
rect 37093 15311 37151 15317
rect 1104 15258 37628 15280
rect 1104 15206 4874 15258
rect 4926 15206 4938 15258
rect 4990 15206 5002 15258
rect 5054 15206 5066 15258
rect 5118 15206 5130 15258
rect 5182 15206 35594 15258
rect 35646 15206 35658 15258
rect 35710 15206 35722 15258
rect 35774 15206 35786 15258
rect 35838 15206 35850 15258
rect 35902 15206 37628 15258
rect 1104 15184 37628 15206
rect 5997 15147 6055 15153
rect 5997 15113 6009 15147
rect 6043 15144 6055 15147
rect 6546 15144 6552 15156
rect 6043 15116 6552 15144
rect 6043 15113 6055 15116
rect 5997 15107 6055 15113
rect 6546 15104 6552 15116
rect 6604 15104 6610 15156
rect 6641 15147 6699 15153
rect 6641 15113 6653 15147
rect 6687 15113 6699 15147
rect 6641 15107 6699 15113
rect 7101 15147 7159 15153
rect 7101 15113 7113 15147
rect 7147 15144 7159 15147
rect 7926 15144 7932 15156
rect 7147 15116 7932 15144
rect 7147 15113 7159 15116
rect 7101 15107 7159 15113
rect 5813 15011 5871 15017
rect 5813 14977 5825 15011
rect 5859 15008 5871 15011
rect 6656 15008 6684 15107
rect 7926 15104 7932 15116
rect 7984 15104 7990 15156
rect 8110 15104 8116 15156
rect 8168 15144 8174 15156
rect 9122 15144 9128 15156
rect 8168 15116 9128 15144
rect 8168 15104 8174 15116
rect 9122 15104 9128 15116
rect 9180 15104 9186 15156
rect 15102 15104 15108 15156
rect 15160 15144 15166 15156
rect 15289 15147 15347 15153
rect 15289 15144 15301 15147
rect 15160 15116 15301 15144
rect 15160 15104 15166 15116
rect 15289 15113 15301 15116
rect 15335 15113 15347 15147
rect 22646 15144 22652 15156
rect 22607 15116 22652 15144
rect 15289 15107 15347 15113
rect 22646 15104 22652 15116
rect 22704 15104 22710 15156
rect 27062 15104 27068 15156
rect 27120 15144 27126 15156
rect 28353 15147 28411 15153
rect 28353 15144 28365 15147
rect 27120 15116 28365 15144
rect 27120 15104 27126 15116
rect 28353 15113 28365 15116
rect 28399 15113 28411 15147
rect 28353 15107 28411 15113
rect 29181 15147 29239 15153
rect 29181 15113 29193 15147
rect 29227 15144 29239 15147
rect 29546 15144 29552 15156
rect 29227 15116 29552 15144
rect 29227 15113 29239 15116
rect 29181 15107 29239 15113
rect 29546 15104 29552 15116
rect 29604 15104 29610 15156
rect 30466 15104 30472 15156
rect 30524 15144 30530 15156
rect 31113 15147 31171 15153
rect 31113 15144 31125 15147
rect 30524 15116 31125 15144
rect 30524 15104 30530 15116
rect 31113 15113 31125 15116
rect 31159 15113 31171 15147
rect 31113 15107 31171 15113
rect 32477 15147 32535 15153
rect 32477 15113 32489 15147
rect 32523 15144 32535 15147
rect 32582 15144 32588 15156
rect 32523 15116 32588 15144
rect 32523 15113 32535 15116
rect 32477 15107 32535 15113
rect 32582 15104 32588 15116
rect 32640 15104 32646 15156
rect 33042 15104 33048 15156
rect 33100 15144 33106 15156
rect 33229 15147 33287 15153
rect 33229 15144 33241 15147
rect 33100 15116 33241 15144
rect 33100 15104 33106 15116
rect 33229 15113 33241 15116
rect 33275 15113 33287 15147
rect 33229 15107 33287 15113
rect 34330 15104 34336 15156
rect 34388 15104 34394 15156
rect 13354 15076 13360 15088
rect 13315 15048 13360 15076
rect 13354 15036 13360 15048
rect 13412 15036 13418 15088
rect 13725 15079 13783 15085
rect 13725 15045 13737 15079
rect 13771 15076 13783 15079
rect 13814 15076 13820 15088
rect 13771 15048 13820 15076
rect 13771 15045 13783 15048
rect 13725 15039 13783 15045
rect 13814 15036 13820 15048
rect 13872 15036 13878 15088
rect 14458 15076 14464 15088
rect 14419 15048 14464 15076
rect 14458 15036 14464 15048
rect 14516 15036 14522 15088
rect 16298 15076 16304 15088
rect 14660 15048 16304 15076
rect 7006 15008 7012 15020
rect 5859 14980 6684 15008
rect 6967 14980 7012 15008
rect 5859 14977 5871 14980
rect 5813 14971 5871 14977
rect 7006 14968 7012 14980
rect 7064 14968 7070 15020
rect 8297 15011 8355 15017
rect 8297 14977 8309 15011
rect 8343 15008 8355 15011
rect 8386 15008 8392 15020
rect 8343 14980 8392 15008
rect 8343 14977 8355 14980
rect 8297 14971 8355 14977
rect 8386 14968 8392 14980
rect 8444 14968 8450 15020
rect 8938 15008 8944 15020
rect 8899 14980 8944 15008
rect 8938 14968 8944 14980
rect 8996 14968 9002 15020
rect 10318 14968 10324 15020
rect 10376 14968 10382 15020
rect 11698 15008 11704 15020
rect 11659 14980 11704 15008
rect 11698 14968 11704 14980
rect 11756 14968 11762 15020
rect 12713 15011 12771 15017
rect 12713 14977 12725 15011
rect 12759 15008 12771 15011
rect 14660 15008 14688 15048
rect 16298 15036 16304 15048
rect 16356 15036 16362 15088
rect 19978 15036 19984 15088
rect 20036 15076 20042 15088
rect 23201 15079 23259 15085
rect 23201 15076 23213 15079
rect 20036 15048 23213 15076
rect 20036 15036 20042 15048
rect 23201 15045 23213 15048
rect 23247 15076 23259 15079
rect 25685 15079 25743 15085
rect 25685 15076 25697 15079
rect 23247 15048 25697 15076
rect 23247 15045 23259 15048
rect 23201 15039 23259 15045
rect 25685 15045 25697 15048
rect 25731 15076 25743 15079
rect 26418 15076 26424 15088
rect 25731 15048 26424 15076
rect 25731 15045 25743 15048
rect 25685 15039 25743 15045
rect 26418 15036 26424 15048
rect 26476 15036 26482 15088
rect 26510 15036 26516 15088
rect 26568 15076 26574 15088
rect 27338 15076 27344 15088
rect 26568 15048 27344 15076
rect 26568 15036 26574 15048
rect 27338 15036 27344 15048
rect 27396 15036 27402 15088
rect 30006 15076 30012 15088
rect 29564 15048 30012 15076
rect 12759 14980 14688 15008
rect 12759 14977 12771 14980
rect 12713 14971 12771 14977
rect 14734 14968 14740 15020
rect 14792 15008 14798 15020
rect 15378 15008 15384 15020
rect 14792 14980 15240 15008
rect 15339 14980 15384 15008
rect 14792 14968 14798 14980
rect 7190 14940 7196 14952
rect 7151 14912 7196 14940
rect 7190 14900 7196 14912
rect 7248 14900 7254 14952
rect 9217 14943 9275 14949
rect 9217 14940 9229 14943
rect 8496 14912 9229 14940
rect 8496 14881 8524 14912
rect 9217 14909 9229 14912
rect 9263 14909 9275 14943
rect 9217 14903 9275 14909
rect 9766 14900 9772 14952
rect 9824 14940 9830 14952
rect 10689 14943 10747 14949
rect 10689 14940 10701 14943
rect 9824 14912 10701 14940
rect 9824 14900 9830 14912
rect 10689 14909 10701 14912
rect 10735 14909 10747 14943
rect 15212 14940 15240 14980
rect 15378 14968 15384 14980
rect 15436 14968 15442 15020
rect 22002 14968 22008 15020
rect 22060 15008 22066 15020
rect 22557 15011 22615 15017
rect 22557 15008 22569 15011
rect 22060 14980 22569 15008
rect 22060 14968 22066 14980
rect 22557 14977 22569 14980
rect 22603 14977 22615 15011
rect 24578 15008 24584 15020
rect 24539 14980 24584 15008
rect 22557 14971 22615 14977
rect 24578 14968 24584 14980
rect 24636 14968 24642 15020
rect 26694 14968 26700 15020
rect 26752 15008 26758 15020
rect 27525 15011 27583 15017
rect 27525 15008 27537 15011
rect 26752 14980 27537 15008
rect 26752 14968 26758 14980
rect 27525 14977 27537 14980
rect 27571 15008 27583 15011
rect 28534 15008 28540 15020
rect 27571 14980 27844 15008
rect 28495 14980 28540 15008
rect 27571 14977 27583 14980
rect 27525 14971 27583 14977
rect 15838 14940 15844 14952
rect 15212 14912 15844 14940
rect 10689 14903 10747 14909
rect 15838 14900 15844 14912
rect 15896 14900 15902 14952
rect 22922 14900 22928 14952
rect 22980 14940 22986 14952
rect 23937 14943 23995 14949
rect 23937 14940 23949 14943
rect 22980 14912 23949 14940
rect 22980 14900 22986 14912
rect 23937 14909 23949 14912
rect 23983 14909 23995 14943
rect 23937 14903 23995 14909
rect 24026 14900 24032 14952
rect 24084 14940 24090 14952
rect 27617 14943 27675 14949
rect 27617 14940 27629 14943
rect 24084 14912 27629 14940
rect 24084 14900 24090 14912
rect 27617 14909 27629 14912
rect 27663 14909 27675 14943
rect 27617 14903 27675 14909
rect 27709 14943 27767 14949
rect 27709 14909 27721 14943
rect 27755 14909 27767 14943
rect 27816 14940 27844 14980
rect 28534 14968 28540 14980
rect 28592 14968 28598 15020
rect 28902 14968 28908 15020
rect 28960 15008 28966 15020
rect 29319 15011 29377 15017
rect 29319 15008 29331 15011
rect 28960 14980 29331 15008
rect 28960 14968 28966 14980
rect 29319 14977 29331 14980
rect 29365 14977 29377 15011
rect 29454 15008 29460 15020
rect 29415 14980 29460 15008
rect 29319 14971 29377 14977
rect 29454 14968 29460 14980
rect 29512 14968 29518 15020
rect 29564 15017 29592 15048
rect 30006 15036 30012 15048
rect 30064 15076 30070 15088
rect 31665 15079 31723 15085
rect 31665 15076 31677 15079
rect 30064 15048 31677 15076
rect 30064 15036 30070 15048
rect 31665 15045 31677 15048
rect 31711 15045 31723 15079
rect 31665 15039 31723 15045
rect 32122 15036 32128 15088
rect 32180 15076 32186 15088
rect 32677 15079 32735 15085
rect 32677 15076 32689 15079
rect 32180 15048 32689 15076
rect 32180 15036 32186 15048
rect 32677 15045 32689 15048
rect 32723 15076 32735 15079
rect 32766 15076 32772 15088
rect 32723 15048 32772 15076
rect 32723 15045 32735 15048
rect 32677 15039 32735 15045
rect 32766 15036 32772 15048
rect 32824 15036 32830 15088
rect 34348 15076 34376 15104
rect 36078 15076 36084 15088
rect 33888 15048 34376 15076
rect 35374 15048 36084 15076
rect 29549 15011 29607 15017
rect 29549 14977 29561 15011
rect 29595 14977 29607 15011
rect 29677 15011 29735 15017
rect 29677 15008 29689 15011
rect 29549 14971 29607 14977
rect 29656 14977 29689 15008
rect 29723 14977 29735 15011
rect 29656 14971 29735 14977
rect 29656 14940 29684 14971
rect 29822 14968 29828 15020
rect 29880 15008 29886 15020
rect 30926 15008 30932 15020
rect 29880 14980 29925 15008
rect 30887 14980 30932 15008
rect 29880 14968 29886 14980
rect 30926 14968 30932 14980
rect 30984 14968 30990 15020
rect 31757 15011 31815 15017
rect 31757 14977 31769 15011
rect 31803 15008 31815 15011
rect 33318 15008 33324 15020
rect 31803 14980 32536 15008
rect 33279 14980 33324 15008
rect 31803 14977 31815 14980
rect 31757 14971 31815 14977
rect 29914 14940 29920 14952
rect 27816 14912 29920 14940
rect 27709 14903 27767 14909
rect 8481 14875 8539 14881
rect 8481 14841 8493 14875
rect 8527 14841 8539 14875
rect 8481 14835 8539 14841
rect 26326 14832 26332 14884
rect 26384 14872 26390 14884
rect 27724 14872 27752 14903
rect 29914 14900 29920 14912
rect 29972 14900 29978 14952
rect 30745 14943 30803 14949
rect 30745 14909 30757 14943
rect 30791 14940 30803 14943
rect 30834 14940 30840 14952
rect 30791 14912 30840 14940
rect 30791 14909 30803 14912
rect 30745 14903 30803 14909
rect 26384 14844 27752 14872
rect 26384 14832 26390 14844
rect 28258 14832 28264 14884
rect 28316 14872 28322 14884
rect 30760 14872 30788 14903
rect 30834 14900 30840 14912
rect 30892 14900 30898 14952
rect 28316 14844 30788 14872
rect 30944 14872 30972 14968
rect 32508 14952 32536 14980
rect 33318 14968 33324 14980
rect 33376 14968 33382 15020
rect 33888 15017 33916 15048
rect 36078 15036 36084 15048
rect 36136 15036 36142 15088
rect 33873 15011 33931 15017
rect 33873 14977 33885 15011
rect 33919 14977 33931 15011
rect 36262 15008 36268 15020
rect 36223 14980 36268 15008
rect 33873 14971 33931 14977
rect 36262 14968 36268 14980
rect 36320 14968 36326 15020
rect 32490 14900 32496 14952
rect 32548 14900 32554 14952
rect 34149 14943 34207 14949
rect 34149 14909 34161 14943
rect 34195 14940 34207 14943
rect 34238 14940 34244 14952
rect 34195 14912 34244 14940
rect 34195 14909 34207 14912
rect 34149 14903 34207 14909
rect 34238 14900 34244 14912
rect 34296 14900 34302 14952
rect 31570 14872 31576 14884
rect 30944 14844 31576 14872
rect 28316 14832 28322 14844
rect 31570 14832 31576 14844
rect 31628 14872 31634 14884
rect 32309 14875 32367 14881
rect 32309 14872 32321 14875
rect 31628 14844 32321 14872
rect 31628 14832 31634 14844
rect 32309 14841 32321 14844
rect 32355 14841 32367 14875
rect 32309 14835 32367 14841
rect 11882 14804 11888 14816
rect 11843 14776 11888 14804
rect 11882 14764 11888 14776
rect 11940 14764 11946 14816
rect 12250 14764 12256 14816
rect 12308 14804 12314 14816
rect 12437 14807 12495 14813
rect 12437 14804 12449 14807
rect 12308 14776 12449 14804
rect 12308 14764 12314 14776
rect 12437 14773 12449 14776
rect 12483 14773 12495 14807
rect 24762 14804 24768 14816
rect 24723 14776 24768 14804
rect 12437 14767 12495 14773
rect 24762 14764 24768 14776
rect 24820 14764 24826 14816
rect 24946 14764 24952 14816
rect 25004 14804 25010 14816
rect 27157 14807 27215 14813
rect 27157 14804 27169 14807
rect 25004 14776 27169 14804
rect 25004 14764 25010 14776
rect 27157 14773 27169 14776
rect 27203 14773 27215 14807
rect 27157 14767 27215 14773
rect 31202 14764 31208 14816
rect 31260 14804 31266 14816
rect 32122 14804 32128 14816
rect 31260 14776 32128 14804
rect 31260 14764 31266 14776
rect 32122 14764 32128 14776
rect 32180 14764 32186 14816
rect 32490 14804 32496 14816
rect 32451 14776 32496 14804
rect 32490 14764 32496 14776
rect 32548 14764 32554 14816
rect 35618 14804 35624 14816
rect 35579 14776 35624 14804
rect 35618 14764 35624 14776
rect 35676 14764 35682 14816
rect 36170 14804 36176 14816
rect 36131 14776 36176 14804
rect 36170 14764 36176 14776
rect 36228 14764 36234 14816
rect 1104 14714 37628 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 37628 14714
rect 1104 14640 37628 14662
rect 6914 14560 6920 14612
rect 6972 14600 6978 14612
rect 7466 14600 7472 14612
rect 6972 14572 7472 14600
rect 6972 14560 6978 14572
rect 7466 14560 7472 14572
rect 7524 14600 7530 14612
rect 7837 14603 7895 14609
rect 7837 14600 7849 14603
rect 7524 14572 7849 14600
rect 7524 14560 7530 14572
rect 7837 14569 7849 14572
rect 7883 14569 7895 14603
rect 11698 14600 11704 14612
rect 11659 14572 11704 14600
rect 7837 14563 7895 14569
rect 11698 14560 11704 14572
rect 11756 14560 11762 14612
rect 21177 14603 21235 14609
rect 21177 14569 21189 14603
rect 21223 14600 21235 14603
rect 24026 14600 24032 14612
rect 21223 14572 24032 14600
rect 21223 14569 21235 14572
rect 21177 14563 21235 14569
rect 24026 14560 24032 14572
rect 24084 14560 24090 14612
rect 25590 14560 25596 14612
rect 25648 14600 25654 14612
rect 27706 14600 27712 14612
rect 25648 14572 27384 14600
rect 27667 14572 27712 14600
rect 25648 14560 25654 14572
rect 2130 14492 2136 14544
rect 2188 14532 2194 14544
rect 10962 14532 10968 14544
rect 2188 14504 6224 14532
rect 2188 14492 2194 14504
rect 6086 14464 6092 14476
rect 6047 14436 6092 14464
rect 6086 14424 6092 14436
rect 6144 14424 6150 14476
rect 6196 14464 6224 14504
rect 9600 14504 10968 14532
rect 9600 14464 9628 14504
rect 10962 14492 10968 14504
rect 11020 14492 11026 14544
rect 13173 14535 13231 14541
rect 13173 14532 13185 14535
rect 12176 14504 13185 14532
rect 9766 14464 9772 14476
rect 6196 14436 9628 14464
rect 9727 14436 9772 14464
rect 9766 14424 9772 14436
rect 9824 14424 9830 14476
rect 9858 14424 9864 14476
rect 9916 14464 9922 14476
rect 10594 14464 10600 14476
rect 9916 14436 10600 14464
rect 9916 14424 9922 14436
rect 10594 14424 10600 14436
rect 10652 14464 10658 14476
rect 11057 14467 11115 14473
rect 11057 14464 11069 14467
rect 10652 14436 11069 14464
rect 10652 14424 10658 14436
rect 11057 14433 11069 14436
rect 11103 14464 11115 14467
rect 12176 14464 12204 14504
rect 13173 14501 13185 14504
rect 13219 14501 13231 14535
rect 13173 14495 13231 14501
rect 11103 14436 12204 14464
rect 11103 14433 11115 14436
rect 11057 14427 11115 14433
rect 12250 14424 12256 14476
rect 12308 14464 12314 14476
rect 12308 14436 12353 14464
rect 12308 14424 12314 14436
rect 21634 14424 21640 14476
rect 21692 14464 21698 14476
rect 22186 14464 22192 14476
rect 21692 14436 22192 14464
rect 21692 14424 21698 14436
rect 22186 14424 22192 14436
rect 22244 14464 22250 14476
rect 22922 14464 22928 14476
rect 22244 14436 22928 14464
rect 22244 14424 22250 14436
rect 22922 14424 22928 14436
rect 22980 14424 22986 14476
rect 24854 14424 24860 14476
rect 24912 14464 24918 14476
rect 24949 14467 25007 14473
rect 24949 14464 24961 14467
rect 24912 14436 24961 14464
rect 24912 14424 24918 14436
rect 24949 14433 24961 14436
rect 24995 14464 25007 14467
rect 26510 14464 26516 14476
rect 24995 14436 26516 14464
rect 24995 14433 25007 14436
rect 24949 14427 25007 14433
rect 26510 14424 26516 14436
rect 26568 14424 26574 14476
rect 5445 14399 5503 14405
rect 5445 14365 5457 14399
rect 5491 14396 5503 14399
rect 5534 14396 5540 14408
rect 5491 14368 5540 14396
rect 5491 14365 5503 14368
rect 5445 14359 5503 14365
rect 5534 14356 5540 14368
rect 5592 14356 5598 14408
rect 8386 14396 8392 14408
rect 8347 14368 8392 14396
rect 8386 14356 8392 14368
rect 8444 14356 8450 14408
rect 10873 14399 10931 14405
rect 10873 14365 10885 14399
rect 10919 14396 10931 14399
rect 11238 14396 11244 14408
rect 10919 14368 11244 14396
rect 10919 14365 10931 14368
rect 10873 14359 10931 14365
rect 11238 14356 11244 14368
rect 11296 14356 11302 14408
rect 13449 14399 13507 14405
rect 13449 14365 13461 14399
rect 13495 14396 13507 14399
rect 13814 14396 13820 14408
rect 13495 14368 13820 14396
rect 13495 14365 13507 14368
rect 13449 14359 13507 14365
rect 13814 14356 13820 14368
rect 13872 14356 13878 14408
rect 21542 14356 21548 14408
rect 21600 14356 21606 14408
rect 23566 14396 23572 14408
rect 23527 14368 23572 14396
rect 23566 14356 23572 14368
rect 23624 14356 23630 14408
rect 27356 14405 27384 14572
rect 27706 14560 27712 14572
rect 27764 14560 27770 14612
rect 28169 14603 28227 14609
rect 28169 14569 28181 14603
rect 28215 14600 28227 14603
rect 28442 14600 28448 14612
rect 28215 14572 28448 14600
rect 28215 14569 28227 14572
rect 28169 14563 28227 14569
rect 28442 14560 28448 14572
rect 28500 14560 28506 14612
rect 28626 14600 28632 14612
rect 28587 14572 28632 14600
rect 28626 14560 28632 14572
rect 28684 14560 28690 14612
rect 31573 14603 31631 14609
rect 31573 14569 31585 14603
rect 31619 14600 31631 14603
rect 31754 14600 31760 14612
rect 31619 14572 31760 14600
rect 31619 14569 31631 14572
rect 31573 14563 31631 14569
rect 31754 14560 31760 14572
rect 31812 14560 31818 14612
rect 32401 14603 32459 14609
rect 32401 14569 32413 14603
rect 32447 14600 32459 14603
rect 34054 14600 34060 14612
rect 32447 14572 34060 14600
rect 32447 14569 32459 14572
rect 32401 14563 32459 14569
rect 34054 14560 34060 14572
rect 34112 14560 34118 14612
rect 34238 14600 34244 14612
rect 34199 14572 34244 14600
rect 34238 14560 34244 14572
rect 34296 14560 34302 14612
rect 35434 14560 35440 14612
rect 35492 14600 35498 14612
rect 35529 14603 35587 14609
rect 35529 14600 35541 14603
rect 35492 14572 35541 14600
rect 35492 14560 35498 14572
rect 35529 14569 35541 14572
rect 35575 14569 35587 14603
rect 35529 14563 35587 14569
rect 28718 14532 28724 14544
rect 28368 14504 28724 14532
rect 27433 14467 27491 14473
rect 27433 14433 27445 14467
rect 27479 14464 27491 14467
rect 28258 14464 28264 14476
rect 27479 14436 28264 14464
rect 27479 14433 27491 14436
rect 27433 14427 27491 14433
rect 28258 14424 28264 14436
rect 28316 14424 28322 14476
rect 28368 14405 28396 14504
rect 28718 14492 28724 14504
rect 28776 14532 28782 14544
rect 31202 14532 31208 14544
rect 28776 14504 31208 14532
rect 28776 14492 28782 14504
rect 31202 14492 31208 14504
rect 31260 14492 31266 14544
rect 34514 14532 34520 14544
rect 31496 14504 34520 14532
rect 29914 14464 29920 14476
rect 29875 14436 29920 14464
rect 29914 14424 29920 14436
rect 29972 14424 29978 14476
rect 30282 14424 30288 14476
rect 30340 14464 30346 14476
rect 30377 14467 30435 14473
rect 30377 14464 30389 14467
rect 30340 14436 30389 14464
rect 30340 14424 30346 14436
rect 30377 14433 30389 14436
rect 30423 14433 30435 14467
rect 30377 14427 30435 14433
rect 27341 14399 27399 14405
rect 27341 14365 27353 14399
rect 27387 14365 27399 14399
rect 27341 14359 27399 14365
rect 28353 14399 28411 14405
rect 28353 14365 28365 14399
rect 28399 14365 28411 14399
rect 28353 14359 28411 14365
rect 28445 14399 28503 14405
rect 28445 14365 28457 14399
rect 28491 14365 28503 14399
rect 28445 14359 28503 14365
rect 28721 14399 28779 14405
rect 28721 14365 28733 14399
rect 28767 14396 28779 14399
rect 28810 14396 28816 14408
rect 28767 14368 28816 14396
rect 28767 14365 28779 14368
rect 28721 14359 28779 14365
rect 6365 14331 6423 14337
rect 6365 14328 6377 14331
rect 5644 14300 6377 14328
rect 5644 14269 5672 14300
rect 6365 14297 6377 14300
rect 6411 14297 6423 14331
rect 6365 14291 6423 14297
rect 7374 14288 7380 14340
rect 7432 14288 7438 14340
rect 9677 14331 9735 14337
rect 9677 14297 9689 14331
rect 9723 14328 9735 14331
rect 10686 14328 10692 14340
rect 9723 14300 10692 14328
rect 9723 14297 9735 14300
rect 9677 14291 9735 14297
rect 10686 14288 10692 14300
rect 10744 14288 10750 14340
rect 12158 14328 12164 14340
rect 12119 14300 12164 14328
rect 12158 14288 12164 14300
rect 12216 14288 12222 14340
rect 22649 14331 22707 14337
rect 22649 14297 22661 14331
rect 22695 14297 22707 14331
rect 25222 14328 25228 14340
rect 25183 14300 25228 14328
rect 22649 14291 22707 14297
rect 5629 14263 5687 14269
rect 5629 14229 5641 14263
rect 5675 14229 5687 14263
rect 8570 14260 8576 14272
rect 8531 14232 8576 14260
rect 5629 14223 5687 14229
rect 8570 14220 8576 14232
rect 8628 14220 8634 14272
rect 9306 14260 9312 14272
rect 9267 14232 9312 14260
rect 9306 14220 9312 14232
rect 9364 14220 9370 14272
rect 10505 14263 10563 14269
rect 10505 14229 10517 14263
rect 10551 14260 10563 14263
rect 10778 14260 10784 14272
rect 10551 14232 10784 14260
rect 10551 14229 10563 14232
rect 10505 14223 10563 14229
rect 10778 14220 10784 14232
rect 10836 14220 10842 14272
rect 10962 14260 10968 14272
rect 10923 14232 10968 14260
rect 10962 14220 10968 14232
rect 11020 14260 11026 14272
rect 12069 14263 12127 14269
rect 12069 14260 12081 14263
rect 11020 14232 12081 14260
rect 11020 14220 11026 14232
rect 12069 14229 12081 14232
rect 12115 14260 12127 14263
rect 13814 14260 13820 14272
rect 12115 14232 13820 14260
rect 12115 14229 12127 14232
rect 12069 14223 12127 14229
rect 13814 14220 13820 14232
rect 13872 14220 13878 14272
rect 22664 14260 22692 14291
rect 25222 14288 25228 14300
rect 25280 14288 25286 14340
rect 27246 14328 27252 14340
rect 26450 14300 27252 14328
rect 27246 14288 27252 14300
rect 27304 14288 27310 14340
rect 28258 14288 28264 14340
rect 28316 14328 28322 14340
rect 28460 14328 28488 14359
rect 28810 14356 28816 14368
rect 28868 14356 28874 14408
rect 29730 14356 29736 14408
rect 29788 14356 29794 14408
rect 30006 14356 30012 14408
rect 30064 14396 30070 14408
rect 31021 14399 31079 14405
rect 30064 14368 30109 14396
rect 30064 14356 30070 14368
rect 31021 14365 31033 14399
rect 31067 14396 31079 14399
rect 31386 14396 31392 14408
rect 31067 14368 31392 14396
rect 31067 14365 31079 14368
rect 31021 14359 31079 14365
rect 31386 14356 31392 14368
rect 31444 14356 31450 14408
rect 28316 14300 28488 14328
rect 29748 14328 29776 14356
rect 30285 14331 30343 14337
rect 30285 14328 30297 14331
rect 29748 14300 30297 14328
rect 28316 14288 28322 14300
rect 30285 14297 30297 14300
rect 30331 14328 30343 14331
rect 31496 14328 31524 14504
rect 34514 14492 34520 14504
rect 34572 14532 34578 14544
rect 35618 14532 35624 14544
rect 34572 14504 35624 14532
rect 34572 14492 34578 14504
rect 35618 14492 35624 14504
rect 35676 14492 35682 14544
rect 31570 14424 31576 14476
rect 31628 14464 31634 14476
rect 31628 14436 32260 14464
rect 31628 14424 31634 14436
rect 32232 14405 32260 14436
rect 32674 14424 32680 14476
rect 32732 14464 32738 14476
rect 34790 14464 34796 14476
rect 32732 14436 34796 14464
rect 32732 14424 32738 14436
rect 31665 14399 31723 14405
rect 31665 14365 31677 14399
rect 31711 14365 31723 14399
rect 31665 14359 31723 14365
rect 32217 14399 32275 14405
rect 32217 14365 32229 14399
rect 32263 14365 32275 14399
rect 32398 14396 32404 14408
rect 32359 14368 32404 14396
rect 32217 14359 32275 14365
rect 30331 14300 31524 14328
rect 31680 14328 31708 14359
rect 32398 14356 32404 14368
rect 32456 14356 32462 14408
rect 32861 14399 32919 14405
rect 32861 14365 32873 14399
rect 32907 14396 32919 14399
rect 33226 14396 33232 14408
rect 32907 14368 33232 14396
rect 32907 14365 32919 14368
rect 32861 14359 32919 14365
rect 33226 14356 33232 14368
rect 33284 14356 33290 14408
rect 34072 14405 34100 14436
rect 34790 14424 34796 14436
rect 34848 14464 34854 14476
rect 35161 14467 35219 14473
rect 35161 14464 35173 14467
rect 34848 14436 35173 14464
rect 34848 14424 34854 14436
rect 35161 14433 35173 14436
rect 35207 14433 35219 14467
rect 35161 14427 35219 14433
rect 34057 14399 34115 14405
rect 34057 14365 34069 14399
rect 34103 14365 34115 14399
rect 34057 14359 34115 14365
rect 34241 14399 34299 14405
rect 34241 14365 34253 14399
rect 34287 14396 34299 14399
rect 34606 14396 34612 14408
rect 34287 14368 34612 14396
rect 34287 14365 34299 14368
rect 34241 14359 34299 14365
rect 34606 14356 34612 14368
rect 34664 14356 34670 14408
rect 35253 14399 35311 14405
rect 35253 14365 35265 14399
rect 35299 14396 35311 14399
rect 36170 14396 36176 14408
rect 35299 14368 36176 14396
rect 35299 14365 35311 14368
rect 35253 14359 35311 14365
rect 36170 14356 36176 14368
rect 36228 14356 36234 14408
rect 33318 14328 33324 14340
rect 31680 14300 33324 14328
rect 30331 14297 30343 14300
rect 30285 14291 30343 14297
rect 33318 14288 33324 14300
rect 33376 14288 33382 14340
rect 23385 14263 23443 14269
rect 23385 14260 23397 14263
rect 22664 14232 23397 14260
rect 23385 14229 23397 14232
rect 23431 14229 23443 14263
rect 26694 14260 26700 14272
rect 26655 14232 26700 14260
rect 23385 14223 23443 14229
rect 26694 14220 26700 14232
rect 26752 14220 26758 14272
rect 29086 14220 29092 14272
rect 29144 14260 29150 14272
rect 29733 14263 29791 14269
rect 29733 14260 29745 14263
rect 29144 14232 29745 14260
rect 29144 14220 29150 14232
rect 29733 14229 29745 14232
rect 29779 14229 29791 14263
rect 29733 14223 29791 14229
rect 30929 14263 30987 14269
rect 30929 14229 30941 14263
rect 30975 14260 30987 14263
rect 31018 14260 31024 14272
rect 30975 14232 31024 14260
rect 30975 14229 30987 14232
rect 30929 14223 30987 14229
rect 31018 14220 31024 14232
rect 31076 14220 31082 14272
rect 33042 14260 33048 14272
rect 33003 14232 33048 14260
rect 33042 14220 33048 14232
rect 33100 14220 33106 14272
rect 1104 14170 37628 14192
rect 1104 14118 4874 14170
rect 4926 14118 4938 14170
rect 4990 14118 5002 14170
rect 5054 14118 5066 14170
rect 5118 14118 5130 14170
rect 5182 14118 35594 14170
rect 35646 14118 35658 14170
rect 35710 14118 35722 14170
rect 35774 14118 35786 14170
rect 35838 14118 35850 14170
rect 35902 14118 37628 14170
rect 1104 14096 37628 14118
rect 7006 14056 7012 14068
rect 6967 14028 7012 14056
rect 7006 14016 7012 14028
rect 7064 14016 7070 14068
rect 7466 14056 7472 14068
rect 7427 14028 7472 14056
rect 7466 14016 7472 14028
rect 7524 14016 7530 14068
rect 8294 14016 8300 14068
rect 8352 14056 8358 14068
rect 9582 14056 9588 14068
rect 8352 14028 9588 14056
rect 8352 14016 8358 14028
rect 9582 14016 9588 14028
rect 9640 14016 9646 14068
rect 10042 14056 10048 14068
rect 10003 14028 10048 14056
rect 10042 14016 10048 14028
rect 10100 14016 10106 14068
rect 10686 14016 10692 14068
rect 10744 14056 10750 14068
rect 11054 14056 11060 14068
rect 10744 14028 11060 14056
rect 10744 14016 10750 14028
rect 11054 14016 11060 14028
rect 11112 14056 11118 14068
rect 12158 14056 12164 14068
rect 11112 14028 12164 14056
rect 11112 14016 11118 14028
rect 12158 14016 12164 14028
rect 12216 14016 12222 14068
rect 13814 14056 13820 14068
rect 13775 14028 13820 14056
rect 13814 14016 13820 14028
rect 13872 14016 13878 14068
rect 21361 14059 21419 14065
rect 21361 14025 21373 14059
rect 21407 14056 21419 14059
rect 21542 14056 21548 14068
rect 21407 14028 21548 14056
rect 21407 14025 21419 14028
rect 21361 14019 21419 14025
rect 21542 14016 21548 14028
rect 21600 14016 21606 14068
rect 22465 14059 22523 14065
rect 22465 14025 22477 14059
rect 22511 14056 22523 14059
rect 23293 14059 23351 14065
rect 23293 14056 23305 14059
rect 22511 14028 23305 14056
rect 22511 14025 22523 14028
rect 22465 14019 22523 14025
rect 23293 14025 23305 14028
rect 23339 14025 23351 14059
rect 23293 14019 23351 14025
rect 23474 14016 23480 14068
rect 23532 14056 23538 14068
rect 23661 14059 23719 14065
rect 23661 14056 23673 14059
rect 23532 14028 23673 14056
rect 23532 14016 23538 14028
rect 23661 14025 23673 14028
rect 23707 14025 23719 14059
rect 23661 14019 23719 14025
rect 23753 14059 23811 14065
rect 23753 14025 23765 14059
rect 23799 14056 23811 14059
rect 26694 14056 26700 14068
rect 23799 14028 26700 14056
rect 23799 14025 23811 14028
rect 23753 14019 23811 14025
rect 26694 14016 26700 14028
rect 26752 14016 26758 14068
rect 27154 14016 27160 14068
rect 27212 14056 27218 14068
rect 30282 14056 30288 14068
rect 27212 14028 29776 14056
rect 30243 14028 30288 14056
rect 27212 14016 27218 14028
rect 8570 13988 8576 14000
rect 8531 13960 8576 13988
rect 8570 13948 8576 13960
rect 8628 13948 8634 14000
rect 9030 13948 9036 14000
rect 9088 13948 9094 14000
rect 11882 13948 11888 14000
rect 11940 13988 11946 14000
rect 12345 13991 12403 13997
rect 12345 13988 12357 13991
rect 11940 13960 12357 13988
rect 11940 13948 11946 13960
rect 12345 13957 12357 13960
rect 12391 13957 12403 13991
rect 13722 13988 13728 14000
rect 13570 13960 13728 13988
rect 12345 13951 12403 13957
rect 13722 13948 13728 13960
rect 13780 13948 13786 14000
rect 22373 13991 22431 13997
rect 22373 13957 22385 13991
rect 22419 13988 22431 13991
rect 24026 13988 24032 14000
rect 22419 13960 24032 13988
rect 22419 13957 22431 13960
rect 22373 13951 22431 13957
rect 24026 13948 24032 13960
rect 24084 13948 24090 14000
rect 24762 13948 24768 14000
rect 24820 13988 24826 14000
rect 25133 13991 25191 13997
rect 25133 13988 25145 13991
rect 24820 13960 25145 13988
rect 24820 13948 24826 13960
rect 25133 13957 25145 13960
rect 25179 13957 25191 13991
rect 29641 13991 29699 13997
rect 29641 13988 29653 13991
rect 26358 13960 29653 13988
rect 25133 13951 25191 13957
rect 29641 13957 29653 13960
rect 29687 13957 29699 13991
rect 29641 13951 29699 13957
rect 7006 13880 7012 13932
rect 7064 13920 7070 13932
rect 7377 13923 7435 13929
rect 7377 13920 7389 13923
rect 7064 13892 7389 13920
rect 7064 13880 7070 13892
rect 7377 13889 7389 13892
rect 7423 13889 7435 13923
rect 8294 13920 8300 13932
rect 8255 13892 8300 13920
rect 7377 13883 7435 13889
rect 8294 13880 8300 13892
rect 8352 13880 8358 13932
rect 10502 13920 10508 13932
rect 10463 13892 10508 13920
rect 10502 13880 10508 13892
rect 10560 13880 10566 13932
rect 13630 13880 13636 13932
rect 13688 13920 13694 13932
rect 14277 13923 14335 13929
rect 14277 13920 14289 13923
rect 13688 13892 14289 13920
rect 13688 13880 13694 13892
rect 14277 13889 14289 13892
rect 14323 13889 14335 13923
rect 14277 13883 14335 13889
rect 21453 13923 21511 13929
rect 21453 13889 21465 13923
rect 21499 13920 21511 13923
rect 22002 13920 22008 13932
rect 21499 13892 22008 13920
rect 21499 13889 21511 13892
rect 21453 13883 21511 13889
rect 22002 13880 22008 13892
rect 22060 13880 22066 13932
rect 24854 13920 24860 13932
rect 24815 13892 24860 13920
rect 24854 13880 24860 13892
rect 24912 13880 24918 13932
rect 26970 13880 26976 13932
rect 27028 13920 27034 13932
rect 27249 13923 27307 13929
rect 27249 13920 27261 13923
rect 27028 13892 27261 13920
rect 27028 13880 27034 13892
rect 27249 13889 27261 13892
rect 27295 13889 27307 13923
rect 28718 13920 28724 13932
rect 28679 13892 28724 13920
rect 27249 13883 27307 13889
rect 28718 13880 28724 13892
rect 28776 13880 28782 13932
rect 28813 13923 28871 13929
rect 28813 13889 28825 13923
rect 28859 13889 28871 13923
rect 28994 13920 29000 13932
rect 28955 13892 29000 13920
rect 28813 13883 28871 13889
rect 7653 13855 7711 13861
rect 7653 13821 7665 13855
rect 7699 13821 7711 13855
rect 7653 13815 7711 13821
rect 7668 13784 7696 13815
rect 9582 13812 9588 13864
rect 9640 13852 9646 13864
rect 12069 13855 12127 13861
rect 12069 13852 12081 13855
rect 9640 13824 12081 13852
rect 9640 13812 9646 13824
rect 12069 13821 12081 13824
rect 12115 13821 12127 13855
rect 12069 13815 12127 13821
rect 7668 13756 7788 13784
rect 7760 13716 7788 13756
rect 8202 13716 8208 13728
rect 7760 13688 8208 13716
rect 8202 13676 8208 13688
rect 8260 13716 8266 13728
rect 9766 13716 9772 13728
rect 8260 13688 9772 13716
rect 8260 13676 8266 13688
rect 9766 13676 9772 13688
rect 9824 13676 9830 13728
rect 10594 13676 10600 13728
rect 10652 13716 10658 13728
rect 10689 13719 10747 13725
rect 10689 13716 10701 13719
rect 10652 13688 10701 13716
rect 10652 13676 10658 13688
rect 10689 13685 10701 13688
rect 10735 13685 10747 13719
rect 12084 13716 12112 13815
rect 13354 13812 13360 13864
rect 13412 13852 13418 13864
rect 14369 13855 14427 13861
rect 14369 13852 14381 13855
rect 13412 13824 14381 13852
rect 13412 13812 13418 13824
rect 14369 13821 14381 13824
rect 14415 13821 14427 13855
rect 14369 13815 14427 13821
rect 22281 13855 22339 13861
rect 22281 13821 22293 13855
rect 22327 13821 22339 13855
rect 23566 13852 23572 13864
rect 22281 13815 22339 13821
rect 22848 13824 23572 13852
rect 22296 13784 22324 13815
rect 22848 13793 22876 13824
rect 23566 13812 23572 13824
rect 23624 13812 23630 13864
rect 23937 13855 23995 13861
rect 23937 13821 23949 13855
rect 23983 13821 23995 13855
rect 26602 13852 26608 13864
rect 26515 13824 26608 13852
rect 23937 13815 23995 13821
rect 22833 13787 22891 13793
rect 22296 13756 22416 13784
rect 12434 13716 12440 13728
rect 12084 13688 12440 13716
rect 10689 13679 10747 13685
rect 12434 13676 12440 13688
rect 12492 13676 12498 13728
rect 22388 13716 22416 13756
rect 22833 13753 22845 13787
rect 22879 13753 22891 13787
rect 22833 13747 22891 13753
rect 23842 13744 23848 13796
rect 23900 13784 23906 13796
rect 23952 13784 23980 13815
rect 26602 13812 26608 13824
rect 26660 13852 26666 13864
rect 27430 13852 27436 13864
rect 26660 13824 27436 13852
rect 26660 13812 26666 13824
rect 27430 13812 27436 13824
rect 27488 13812 27494 13864
rect 27525 13855 27583 13861
rect 27525 13821 27537 13855
rect 27571 13852 27583 13855
rect 27614 13852 27620 13864
rect 27571 13824 27620 13852
rect 27571 13821 27583 13824
rect 27525 13815 27583 13821
rect 27614 13812 27620 13824
rect 27672 13812 27678 13864
rect 28258 13812 28264 13864
rect 28316 13852 28322 13864
rect 28828 13852 28856 13883
rect 28994 13880 29000 13892
rect 29052 13880 29058 13932
rect 29086 13880 29092 13932
rect 29144 13920 29150 13932
rect 29549 13923 29607 13929
rect 29144 13892 29189 13920
rect 29144 13880 29150 13892
rect 29549 13889 29561 13923
rect 29595 13920 29607 13923
rect 29748 13920 29776 14028
rect 30282 14016 30288 14028
rect 30340 14016 30346 14068
rect 33226 14056 33232 14068
rect 33187 14028 33232 14056
rect 33226 14016 33232 14028
rect 33284 14016 33290 14068
rect 31386 13948 31392 14000
rect 31444 13988 31450 14000
rect 31444 13960 33824 13988
rect 31444 13948 31450 13960
rect 29595 13892 29776 13920
rect 30193 13923 30251 13929
rect 29595 13889 29607 13892
rect 29549 13883 29607 13889
rect 30193 13889 30205 13923
rect 30239 13920 30251 13923
rect 30282 13920 30288 13932
rect 30239 13892 30288 13920
rect 30239 13889 30251 13892
rect 30193 13883 30251 13889
rect 30282 13880 30288 13892
rect 30340 13880 30346 13932
rect 30558 13880 30564 13932
rect 30616 13920 30622 13932
rect 31021 13923 31079 13929
rect 31021 13920 31033 13923
rect 30616 13892 31033 13920
rect 30616 13880 30622 13892
rect 31021 13889 31033 13892
rect 31067 13889 31079 13923
rect 31478 13920 31484 13932
rect 31439 13892 31484 13920
rect 31021 13883 31079 13889
rect 31478 13880 31484 13892
rect 31536 13880 31542 13932
rect 32030 13880 32036 13932
rect 32088 13920 32094 13932
rect 33796 13929 33824 13960
rect 32861 13923 32919 13929
rect 32861 13920 32873 13923
rect 32088 13892 32873 13920
rect 32088 13880 32094 13892
rect 32861 13889 32873 13892
rect 32907 13889 32919 13923
rect 32861 13883 32919 13889
rect 33781 13923 33839 13929
rect 33781 13889 33793 13923
rect 33827 13920 33839 13923
rect 34790 13920 34796 13932
rect 33827 13892 34796 13920
rect 33827 13889 33839 13892
rect 33781 13883 33839 13889
rect 34790 13880 34796 13892
rect 34848 13880 34854 13932
rect 28316 13824 28856 13852
rect 32585 13855 32643 13861
rect 28316 13812 28322 13824
rect 32585 13821 32597 13855
rect 32631 13821 32643 13855
rect 32766 13852 32772 13864
rect 32727 13824 32772 13852
rect 32585 13815 32643 13821
rect 23900 13756 23980 13784
rect 28537 13787 28595 13793
rect 23900 13744 23906 13756
rect 28537 13753 28549 13787
rect 28583 13784 28595 13787
rect 29178 13784 29184 13796
rect 28583 13756 29184 13784
rect 28583 13753 28595 13756
rect 28537 13747 28595 13753
rect 29178 13744 29184 13756
rect 29236 13744 29242 13796
rect 31202 13784 31208 13796
rect 29288 13756 31208 13784
rect 23382 13716 23388 13728
rect 22388 13688 23388 13716
rect 23382 13676 23388 13688
rect 23440 13676 23446 13728
rect 28350 13676 28356 13728
rect 28408 13716 28414 13728
rect 29288 13716 29316 13756
rect 31202 13744 31208 13756
rect 31260 13744 31266 13796
rect 32122 13744 32128 13796
rect 32180 13784 32186 13796
rect 32600 13784 32628 13815
rect 32766 13812 32772 13824
rect 32824 13812 32830 13864
rect 32180 13756 32628 13784
rect 32180 13744 32186 13756
rect 32674 13744 32680 13796
rect 32732 13784 32738 13796
rect 32732 13756 34008 13784
rect 32732 13744 32738 13756
rect 30834 13716 30840 13728
rect 28408 13688 29316 13716
rect 30795 13688 30840 13716
rect 28408 13676 28414 13688
rect 30834 13676 30840 13688
rect 30892 13676 30898 13728
rect 31662 13716 31668 13728
rect 31623 13688 31668 13716
rect 31662 13676 31668 13688
rect 31720 13676 31726 13728
rect 33778 13676 33784 13728
rect 33836 13716 33842 13728
rect 33873 13719 33931 13725
rect 33873 13716 33885 13719
rect 33836 13688 33885 13716
rect 33836 13676 33842 13688
rect 33873 13685 33885 13688
rect 33919 13685 33931 13719
rect 33980 13716 34008 13756
rect 34514 13744 34520 13796
rect 34572 13784 34578 13796
rect 36814 13784 36820 13796
rect 34572 13756 36820 13784
rect 34572 13744 34578 13756
rect 36814 13744 36820 13756
rect 36872 13744 36878 13796
rect 36998 13716 37004 13728
rect 33980 13688 37004 13716
rect 33873 13679 33931 13685
rect 36998 13676 37004 13688
rect 37056 13676 37062 13728
rect 1104 13626 37628 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 37628 13626
rect 1104 13552 37628 13574
rect 7285 13515 7343 13521
rect 7285 13481 7297 13515
rect 7331 13512 7343 13515
rect 7374 13512 7380 13524
rect 7331 13484 7380 13512
rect 7331 13481 7343 13484
rect 7285 13475 7343 13481
rect 7374 13472 7380 13484
rect 7432 13472 7438 13524
rect 8386 13472 8392 13524
rect 8444 13512 8450 13524
rect 9125 13515 9183 13521
rect 9125 13512 9137 13515
rect 8444 13484 9137 13512
rect 8444 13472 8450 13484
rect 9125 13481 9137 13484
rect 9171 13481 9183 13515
rect 9125 13475 9183 13481
rect 9674 13472 9680 13524
rect 9732 13472 9738 13524
rect 12069 13515 12127 13521
rect 12069 13481 12081 13515
rect 12115 13512 12127 13515
rect 12158 13512 12164 13524
rect 12115 13484 12164 13512
rect 12115 13481 12127 13484
rect 12069 13475 12127 13481
rect 12158 13472 12164 13484
rect 12216 13472 12222 13524
rect 24578 13512 24584 13524
rect 24539 13484 24584 13512
rect 24578 13472 24584 13484
rect 24636 13472 24642 13524
rect 26145 13515 26203 13521
rect 26145 13481 26157 13515
rect 26191 13512 26203 13515
rect 26326 13512 26332 13524
rect 26191 13484 26332 13512
rect 26191 13481 26203 13484
rect 26145 13475 26203 13481
rect 2222 13404 2228 13456
rect 2280 13444 2286 13456
rect 8294 13444 8300 13456
rect 2280 13416 8300 13444
rect 2280 13404 2286 13416
rect 8294 13404 8300 13416
rect 8352 13404 8358 13456
rect 8481 13447 8539 13453
rect 8481 13413 8493 13447
rect 8527 13444 8539 13447
rect 9030 13444 9036 13456
rect 8527 13416 9036 13444
rect 8527 13413 8539 13416
rect 8481 13407 8539 13413
rect 9030 13404 9036 13416
rect 9088 13404 9094 13456
rect 9692 13444 9720 13472
rect 22465 13447 22523 13453
rect 22465 13444 22477 13447
rect 9692 13416 10364 13444
rect 10336 13385 10364 13416
rect 22066 13416 22477 13444
rect 9769 13379 9827 13385
rect 9769 13345 9781 13379
rect 9815 13376 9827 13379
rect 10321 13379 10379 13385
rect 9815 13348 10272 13376
rect 9815 13345 9827 13348
rect 9769 13339 9827 13345
rect 1765 13311 1823 13317
rect 1765 13277 1777 13311
rect 1811 13277 1823 13311
rect 1765 13271 1823 13277
rect 1780 13240 1808 13271
rect 5810 13268 5816 13320
rect 5868 13308 5874 13320
rect 6549 13311 6607 13317
rect 6549 13308 6561 13311
rect 5868 13280 6561 13308
rect 5868 13268 5874 13280
rect 6549 13277 6561 13280
rect 6595 13277 6607 13311
rect 6549 13271 6607 13277
rect 7282 13268 7288 13320
rect 7340 13308 7346 13320
rect 7377 13311 7435 13317
rect 7377 13308 7389 13311
rect 7340 13280 7389 13308
rect 7340 13268 7346 13280
rect 7377 13277 7389 13280
rect 7423 13277 7435 13311
rect 8570 13308 8576 13320
rect 8531 13280 8576 13308
rect 7377 13271 7435 13277
rect 8570 13268 8576 13280
rect 8628 13268 8634 13320
rect 9306 13268 9312 13320
rect 9364 13308 9370 13320
rect 9493 13311 9551 13317
rect 9493 13308 9505 13311
rect 9364 13280 9505 13308
rect 9364 13268 9370 13280
rect 9493 13277 9505 13280
rect 9539 13277 9551 13311
rect 9493 13271 9551 13277
rect 9585 13311 9643 13317
rect 9585 13277 9597 13311
rect 9631 13308 9643 13311
rect 10042 13308 10048 13320
rect 9631 13280 10048 13308
rect 9631 13277 9643 13280
rect 9585 13271 9643 13277
rect 10042 13268 10048 13280
rect 10100 13268 10106 13320
rect 8478 13240 8484 13252
rect 1780 13212 8484 13240
rect 8478 13200 8484 13212
rect 8536 13200 8542 13252
rect 10244 13240 10272 13348
rect 10321 13345 10333 13379
rect 10367 13345 10379 13379
rect 10594 13376 10600 13388
rect 10555 13348 10600 13376
rect 10321 13339 10379 13345
rect 10594 13336 10600 13348
rect 10652 13336 10658 13388
rect 12434 13268 12440 13320
rect 12492 13308 12498 13320
rect 13449 13311 13507 13317
rect 13449 13308 13461 13311
rect 12492 13280 13461 13308
rect 12492 13268 12498 13280
rect 13449 13277 13461 13280
rect 13495 13277 13507 13311
rect 13449 13271 13507 13277
rect 13814 13268 13820 13320
rect 13872 13308 13878 13320
rect 14369 13311 14427 13317
rect 14369 13308 14381 13311
rect 13872 13280 14381 13308
rect 13872 13268 13878 13280
rect 14369 13277 14381 13280
rect 14415 13308 14427 13311
rect 14642 13308 14648 13320
rect 14415 13280 14648 13308
rect 14415 13277 14427 13280
rect 14369 13271 14427 13277
rect 14642 13268 14648 13280
rect 14700 13268 14706 13320
rect 21913 13311 21971 13317
rect 21913 13277 21925 13311
rect 21959 13308 21971 13311
rect 22066 13308 22094 13416
rect 22465 13413 22477 13416
rect 22511 13413 22523 13447
rect 22465 13407 22523 13413
rect 24029 13447 24087 13453
rect 24029 13413 24041 13447
rect 24075 13444 24087 13447
rect 25222 13444 25228 13456
rect 24075 13416 25228 13444
rect 24075 13413 24087 13416
rect 24029 13407 24087 13413
rect 25222 13404 25228 13416
rect 25280 13404 25286 13456
rect 23106 13376 23112 13388
rect 23019 13348 23112 13376
rect 23106 13336 23112 13348
rect 23164 13376 23170 13388
rect 23382 13376 23388 13388
rect 23164 13348 23388 13376
rect 23164 13336 23170 13348
rect 23382 13336 23388 13348
rect 23440 13336 23446 13388
rect 25133 13379 25191 13385
rect 25133 13345 25145 13379
rect 25179 13376 25191 13379
rect 26160 13376 26188 13475
rect 26326 13472 26332 13484
rect 26384 13472 26390 13524
rect 27065 13515 27123 13521
rect 27065 13481 27077 13515
rect 27111 13512 27123 13515
rect 27522 13512 27528 13524
rect 27111 13484 27528 13512
rect 27111 13481 27123 13484
rect 27065 13475 27123 13481
rect 27522 13472 27528 13484
rect 27580 13512 27586 13524
rect 28810 13512 28816 13524
rect 27580 13484 28816 13512
rect 27580 13472 27586 13484
rect 28810 13472 28816 13484
rect 28868 13472 28874 13524
rect 30466 13472 30472 13524
rect 30524 13512 30530 13524
rect 31481 13515 31539 13521
rect 31481 13512 31493 13515
rect 30524 13484 31493 13512
rect 30524 13472 30530 13484
rect 31481 13481 31493 13484
rect 31527 13512 31539 13515
rect 32674 13512 32680 13524
rect 31527 13484 32680 13512
rect 31527 13481 31539 13484
rect 31481 13475 31539 13481
rect 32674 13472 32680 13484
rect 32732 13472 32738 13524
rect 32766 13472 32772 13524
rect 32824 13512 32830 13524
rect 33226 13512 33232 13524
rect 32824 13484 33232 13512
rect 32824 13472 32830 13484
rect 33226 13472 33232 13484
rect 33284 13512 33290 13524
rect 33689 13515 33747 13521
rect 33689 13512 33701 13515
rect 33284 13484 33701 13512
rect 33284 13472 33290 13484
rect 33689 13481 33701 13484
rect 33735 13481 33747 13515
rect 33689 13475 33747 13481
rect 31202 13404 31208 13456
rect 31260 13444 31266 13456
rect 31260 13416 32076 13444
rect 31260 13404 31266 13416
rect 25179 13348 26188 13376
rect 25179 13345 25191 13348
rect 25133 13339 25191 13345
rect 27338 13336 27344 13388
rect 27396 13376 27402 13388
rect 28813 13379 28871 13385
rect 28813 13376 28825 13379
rect 27396 13348 28825 13376
rect 27396 13336 27402 13348
rect 28813 13345 28825 13348
rect 28859 13376 28871 13379
rect 29733 13379 29791 13385
rect 29733 13376 29745 13379
rect 28859 13348 29745 13376
rect 28859 13345 28871 13348
rect 28813 13339 28871 13345
rect 29733 13345 29745 13348
rect 29779 13376 29791 13379
rect 32048 13376 32076 13416
rect 29779 13348 31754 13376
rect 32048 13348 34376 13376
rect 29779 13345 29791 13348
rect 29733 13339 29791 13345
rect 21959 13280 22094 13308
rect 23845 13311 23903 13317
rect 21959 13277 21971 13280
rect 21913 13271 21971 13277
rect 23845 13277 23857 13311
rect 23891 13308 23903 13311
rect 24946 13308 24952 13320
rect 23891 13280 24952 13308
rect 23891 13277 23903 13280
rect 23845 13271 23903 13277
rect 24946 13268 24952 13280
rect 25004 13268 25010 13320
rect 26602 13308 26608 13320
rect 25792 13280 26608 13308
rect 10594 13240 10600 13252
rect 10244 13212 10600 13240
rect 10594 13200 10600 13212
rect 10652 13200 10658 13252
rect 11822 13212 12434 13240
rect 1578 13172 1584 13184
rect 1539 13144 1584 13172
rect 1578 13132 1584 13144
rect 1636 13132 1642 13184
rect 6641 13175 6699 13181
rect 6641 13141 6653 13175
rect 6687 13172 6699 13175
rect 7098 13172 7104 13184
rect 6687 13144 7104 13172
rect 6687 13141 6699 13144
rect 6641 13135 6699 13141
rect 7098 13132 7104 13144
rect 7156 13132 7162 13184
rect 12406 13172 12434 13212
rect 12618 13200 12624 13252
rect 12676 13240 12682 13252
rect 12713 13243 12771 13249
rect 12713 13240 12725 13243
rect 12676 13212 12725 13240
rect 12676 13200 12682 13212
rect 12713 13209 12725 13212
rect 12759 13209 12771 13243
rect 25792 13240 25820 13280
rect 26602 13268 26608 13280
rect 26660 13268 26666 13320
rect 31726 13308 31754 13348
rect 34348 13320 34376 13348
rect 31938 13308 31944 13320
rect 31726 13280 31944 13308
rect 31938 13268 31944 13280
rect 31996 13268 32002 13320
rect 34330 13308 34336 13320
rect 34243 13280 34336 13308
rect 34330 13268 34336 13280
rect 34388 13268 34394 13320
rect 34422 13268 34428 13320
rect 34480 13308 34486 13320
rect 36909 13311 36967 13317
rect 36909 13308 36921 13311
rect 34480 13280 36921 13308
rect 34480 13268 34486 13280
rect 36909 13277 36921 13280
rect 36955 13277 36967 13311
rect 36909 13271 36967 13277
rect 12713 13203 12771 13209
rect 24964 13212 25820 13240
rect 13354 13172 13360 13184
rect 12406 13144 13360 13172
rect 13354 13132 13360 13144
rect 13412 13132 13418 13184
rect 14182 13132 14188 13184
rect 14240 13172 14246 13184
rect 14461 13175 14519 13181
rect 14461 13172 14473 13175
rect 14240 13144 14473 13172
rect 14240 13132 14246 13144
rect 14461 13141 14473 13144
rect 14507 13141 14519 13175
rect 14461 13135 14519 13141
rect 21450 13132 21456 13184
rect 21508 13172 21514 13184
rect 21729 13175 21787 13181
rect 21729 13172 21741 13175
rect 21508 13144 21741 13172
rect 21508 13132 21514 13144
rect 21729 13141 21741 13144
rect 21775 13141 21787 13175
rect 22830 13172 22836 13184
rect 22791 13144 22836 13172
rect 21729 13135 21787 13141
rect 22830 13132 22836 13144
rect 22888 13132 22894 13184
rect 22922 13132 22928 13184
rect 22980 13172 22986 13184
rect 22980 13144 23025 13172
rect 22980 13132 22986 13144
rect 23658 13132 23664 13184
rect 23716 13172 23722 13184
rect 24964 13181 24992 13212
rect 25866 13200 25872 13252
rect 25924 13240 25930 13252
rect 25924 13212 25969 13240
rect 25924 13200 25930 13212
rect 26326 13200 26332 13252
rect 26384 13240 26390 13252
rect 26786 13240 26792 13252
rect 26384 13212 26792 13240
rect 26384 13200 26390 13212
rect 26786 13200 26792 13212
rect 26844 13200 26850 13252
rect 28537 13243 28595 13249
rect 28106 13212 28212 13240
rect 24949 13175 25007 13181
rect 24949 13172 24961 13175
rect 23716 13144 24961 13172
rect 23716 13132 23722 13144
rect 24949 13141 24961 13144
rect 24995 13141 25007 13175
rect 24949 13135 25007 13141
rect 25038 13132 25044 13184
rect 25096 13172 25102 13184
rect 28184 13172 28212 13212
rect 28537 13209 28549 13243
rect 28583 13240 28595 13243
rect 28810 13240 28816 13252
rect 28583 13212 28816 13240
rect 28583 13209 28595 13212
rect 28537 13203 28595 13209
rect 28810 13200 28816 13212
rect 28868 13200 28874 13252
rect 30009 13243 30067 13249
rect 30009 13209 30021 13243
rect 30055 13209 30067 13243
rect 30009 13203 30067 13209
rect 29086 13172 29092 13184
rect 25096 13144 25141 13172
rect 28184 13144 29092 13172
rect 25096 13132 25102 13144
rect 29086 13132 29092 13144
rect 29144 13132 29150 13184
rect 30024 13172 30052 13203
rect 31018 13200 31024 13252
rect 31076 13200 31082 13252
rect 31662 13200 31668 13252
rect 31720 13240 31726 13252
rect 32217 13243 32275 13249
rect 32217 13240 32229 13243
rect 31720 13212 32229 13240
rect 31720 13200 31726 13212
rect 32217 13209 32229 13212
rect 32263 13209 32275 13243
rect 34241 13243 34299 13249
rect 34241 13240 34253 13243
rect 33442 13212 34253 13240
rect 32217 13203 32275 13209
rect 34241 13209 34253 13212
rect 34287 13209 34299 13243
rect 34241 13203 34299 13209
rect 30834 13172 30840 13184
rect 30024 13144 30840 13172
rect 30834 13132 30840 13144
rect 30892 13132 30898 13184
rect 37090 13172 37096 13184
rect 37051 13144 37096 13172
rect 37090 13132 37096 13144
rect 37148 13132 37154 13184
rect 1104 13082 37628 13104
rect 1104 13030 4874 13082
rect 4926 13030 4938 13082
rect 4990 13030 5002 13082
rect 5054 13030 5066 13082
rect 5118 13030 5130 13082
rect 5182 13030 35594 13082
rect 35646 13030 35658 13082
rect 35710 13030 35722 13082
rect 35774 13030 35786 13082
rect 35838 13030 35850 13082
rect 35902 13030 37628 13082
rect 1104 13008 37628 13030
rect 9493 12971 9551 12977
rect 9493 12937 9505 12971
rect 9539 12968 9551 12971
rect 10042 12968 10048 12980
rect 9539 12940 10048 12968
rect 9539 12937 9551 12940
rect 9493 12931 9551 12937
rect 10042 12928 10048 12940
rect 10100 12928 10106 12980
rect 10413 12971 10471 12977
rect 10413 12937 10425 12971
rect 10459 12968 10471 12971
rect 10502 12968 10508 12980
rect 10459 12940 10508 12968
rect 10459 12937 10471 12940
rect 10413 12931 10471 12937
rect 10502 12928 10508 12940
rect 10560 12928 10566 12980
rect 10778 12968 10784 12980
rect 10739 12940 10784 12968
rect 10778 12928 10784 12940
rect 10836 12928 10842 12980
rect 10873 12971 10931 12977
rect 10873 12937 10885 12971
rect 10919 12968 10931 12971
rect 11054 12968 11060 12980
rect 10919 12940 11060 12968
rect 10919 12937 10931 12940
rect 10873 12931 10931 12937
rect 11054 12928 11060 12940
rect 11112 12928 11118 12980
rect 13722 12928 13728 12980
rect 13780 12968 13786 12980
rect 14277 12971 14335 12977
rect 14277 12968 14289 12971
rect 13780 12940 14289 12968
rect 13780 12928 13786 12940
rect 14277 12937 14289 12940
rect 14323 12937 14335 12971
rect 14277 12931 14335 12937
rect 22830 12928 22836 12980
rect 22888 12968 22894 12980
rect 23201 12971 23259 12977
rect 23201 12968 23213 12971
rect 22888 12940 23213 12968
rect 22888 12928 22894 12940
rect 23201 12937 23213 12940
rect 23247 12937 23259 12971
rect 23658 12968 23664 12980
rect 23619 12940 23664 12968
rect 23201 12931 23259 12937
rect 23658 12928 23664 12940
rect 23716 12928 23722 12980
rect 25866 12968 25872 12980
rect 25827 12940 25872 12968
rect 25866 12928 25872 12940
rect 25924 12928 25930 12980
rect 27246 12968 27252 12980
rect 27207 12940 27252 12968
rect 27246 12928 27252 12940
rect 27304 12928 27310 12980
rect 28258 12968 28264 12980
rect 28219 12940 28264 12968
rect 28258 12928 28264 12940
rect 28316 12928 28322 12980
rect 28810 12968 28816 12980
rect 28771 12940 28816 12968
rect 28810 12928 28816 12940
rect 28868 12928 28874 12980
rect 30558 12968 30564 12980
rect 30519 12940 30564 12968
rect 30558 12928 30564 12940
rect 30616 12928 30622 12980
rect 31478 12928 31484 12980
rect 31536 12968 31542 12980
rect 31757 12971 31815 12977
rect 31757 12968 31769 12971
rect 31536 12940 31769 12968
rect 31536 12928 31542 12940
rect 31757 12937 31769 12940
rect 31803 12937 31815 12971
rect 33226 12968 33232 12980
rect 31757 12931 31815 12937
rect 32876 12940 33232 12968
rect 7098 12860 7104 12912
rect 7156 12900 7162 12912
rect 7156 12872 7314 12900
rect 7156 12860 7162 12872
rect 8294 12860 8300 12912
rect 8352 12900 8358 12912
rect 12069 12903 12127 12909
rect 12069 12900 12081 12903
rect 8352 12872 12081 12900
rect 8352 12860 8358 12872
rect 12069 12869 12081 12872
rect 12115 12900 12127 12903
rect 12802 12900 12808 12912
rect 12115 12872 12808 12900
rect 12115 12869 12127 12872
rect 12069 12863 12127 12869
rect 12802 12860 12808 12872
rect 12860 12900 12866 12912
rect 13538 12900 13544 12912
rect 12860 12872 13544 12900
rect 12860 12860 12866 12872
rect 13538 12860 13544 12872
rect 13596 12860 13602 12912
rect 22922 12860 22928 12912
rect 22980 12900 22986 12912
rect 24765 12903 24823 12909
rect 24765 12900 24777 12903
rect 22980 12872 24777 12900
rect 22980 12860 22986 12872
rect 24765 12869 24777 12872
rect 24811 12900 24823 12903
rect 25038 12900 25044 12912
rect 24811 12872 25044 12900
rect 24811 12869 24823 12872
rect 24765 12863 24823 12869
rect 25038 12860 25044 12872
rect 25096 12860 25102 12912
rect 31297 12903 31355 12909
rect 31297 12869 31309 12903
rect 31343 12900 31355 12903
rect 32876 12900 32904 12940
rect 33226 12928 33232 12940
rect 33284 12928 33290 12980
rect 34514 12968 34520 12980
rect 34475 12940 34520 12968
rect 34514 12928 34520 12940
rect 34572 12928 34578 12980
rect 33042 12900 33048 12912
rect 31343 12872 32904 12900
rect 33003 12872 33048 12900
rect 31343 12869 31355 12872
rect 31297 12863 31355 12869
rect 33042 12860 33048 12872
rect 33100 12860 33106 12912
rect 33778 12860 33784 12912
rect 33836 12860 33842 12912
rect 6086 12792 6092 12844
rect 6144 12832 6150 12844
rect 6546 12832 6552 12844
rect 6144 12804 6552 12832
rect 6144 12792 6150 12804
rect 6546 12792 6552 12804
rect 6604 12792 6610 12844
rect 11054 12792 11060 12844
rect 11112 12832 11118 12844
rect 12250 12838 12256 12844
rect 12176 12832 12256 12838
rect 11112 12804 12256 12832
rect 11112 12792 11118 12804
rect 12250 12792 12256 12804
rect 12308 12832 12314 12844
rect 12308 12804 12388 12832
rect 12308 12792 12314 12804
rect 6822 12764 6828 12776
rect 6783 12736 6828 12764
rect 6822 12724 6828 12736
rect 6880 12724 6886 12776
rect 8478 12724 8484 12776
rect 8536 12764 8542 12776
rect 9490 12764 9496 12776
rect 8536 12736 9496 12764
rect 8536 12724 8542 12736
rect 9490 12724 9496 12736
rect 9548 12764 9554 12776
rect 9585 12767 9643 12773
rect 9585 12764 9597 12767
rect 9548 12736 9597 12764
rect 9548 12724 9554 12736
rect 9585 12733 9597 12736
rect 9631 12733 9643 12767
rect 9766 12764 9772 12776
rect 9727 12736 9772 12764
rect 9585 12727 9643 12733
rect 9766 12724 9772 12736
rect 9824 12724 9830 12776
rect 10965 12767 11023 12773
rect 10965 12733 10977 12767
rect 11011 12733 11023 12767
rect 10965 12727 11023 12733
rect 10594 12656 10600 12708
rect 10652 12696 10658 12708
rect 10980 12696 11008 12727
rect 11238 12724 11244 12776
rect 11296 12764 11302 12776
rect 12360 12773 12388 12804
rect 13078 12792 13084 12844
rect 13136 12832 13142 12844
rect 13449 12835 13507 12841
rect 13449 12832 13461 12835
rect 13136 12804 13461 12832
rect 13136 12792 13142 12804
rect 13449 12801 13461 12804
rect 13495 12801 13507 12835
rect 13449 12795 13507 12801
rect 13725 12835 13783 12841
rect 13725 12801 13737 12835
rect 13771 12832 13783 12835
rect 13814 12832 13820 12844
rect 13771 12804 13820 12832
rect 13771 12801 13783 12804
rect 13725 12795 13783 12801
rect 13814 12792 13820 12804
rect 13872 12792 13878 12844
rect 14369 12835 14427 12841
rect 14369 12801 14381 12835
rect 14415 12832 14427 12835
rect 14458 12832 14464 12844
rect 14415 12804 14464 12832
rect 14415 12801 14427 12804
rect 14369 12795 14427 12801
rect 14458 12792 14464 12804
rect 14516 12792 14522 12844
rect 14642 12792 14648 12844
rect 14700 12832 14706 12844
rect 17773 12835 17831 12841
rect 17773 12832 17785 12835
rect 14700 12804 17785 12832
rect 14700 12792 14706 12804
rect 17773 12801 17785 12804
rect 17819 12801 17831 12835
rect 17773 12795 17831 12801
rect 22094 12792 22100 12844
rect 22152 12832 22158 12844
rect 22830 12832 22836 12844
rect 22152 12804 22836 12832
rect 22152 12792 22158 12804
rect 22830 12792 22836 12804
rect 22888 12792 22894 12844
rect 23569 12835 23627 12841
rect 23569 12801 23581 12835
rect 23615 12832 23627 12835
rect 24026 12832 24032 12844
rect 23615 12804 24032 12832
rect 23615 12801 23627 12804
rect 23569 12795 23627 12801
rect 24026 12792 24032 12804
rect 24084 12792 24090 12844
rect 24946 12832 24952 12844
rect 24504 12804 24952 12832
rect 12161 12767 12219 12773
rect 12161 12764 12173 12767
rect 11296 12736 12173 12764
rect 11296 12724 11302 12736
rect 12161 12733 12173 12736
rect 12207 12733 12219 12767
rect 12161 12727 12219 12733
rect 12345 12767 12403 12773
rect 12345 12733 12357 12767
rect 12391 12733 12403 12767
rect 12345 12727 12403 12733
rect 17589 12767 17647 12773
rect 17589 12733 17601 12767
rect 17635 12764 17647 12767
rect 18690 12764 18696 12776
rect 17635 12736 18696 12764
rect 17635 12733 17647 12736
rect 17589 12727 17647 12733
rect 18690 12724 18696 12736
rect 18748 12724 18754 12776
rect 23842 12764 23848 12776
rect 23803 12736 23848 12764
rect 23842 12724 23848 12736
rect 23900 12764 23906 12776
rect 24504 12764 24532 12804
rect 24946 12792 24952 12804
rect 25004 12832 25010 12844
rect 25961 12835 26019 12841
rect 25004 12804 25084 12832
rect 25004 12792 25010 12804
rect 23900 12736 24532 12764
rect 23900 12724 23906 12736
rect 24578 12724 24584 12776
rect 24636 12764 24642 12776
rect 25056 12773 25084 12804
rect 25961 12801 25973 12835
rect 26007 12832 26019 12835
rect 26050 12832 26056 12844
rect 26007 12804 26056 12832
rect 26007 12801 26019 12804
rect 25961 12795 26019 12801
rect 26050 12792 26056 12804
rect 26108 12792 26114 12844
rect 27154 12792 27160 12844
rect 27212 12832 27218 12844
rect 27341 12835 27399 12841
rect 27341 12832 27353 12835
rect 27212 12804 27353 12832
rect 27212 12792 27218 12804
rect 27341 12801 27353 12804
rect 27387 12801 27399 12835
rect 27341 12795 27399 12801
rect 27430 12792 27436 12844
rect 27488 12832 27494 12844
rect 28169 12835 28227 12841
rect 28169 12832 28181 12835
rect 27488 12804 28181 12832
rect 27488 12792 27494 12804
rect 28169 12801 28181 12804
rect 28215 12801 28227 12835
rect 28994 12832 29000 12844
rect 28955 12804 29000 12832
rect 28169 12795 28227 12801
rect 28994 12792 29000 12804
rect 29052 12792 29058 12844
rect 30193 12835 30251 12841
rect 30193 12801 30205 12835
rect 30239 12832 30251 12835
rect 30466 12832 30472 12844
rect 30239 12804 30472 12832
rect 30239 12801 30251 12804
rect 30193 12795 30251 12801
rect 30466 12792 30472 12804
rect 30524 12792 30530 12844
rect 31386 12832 31392 12844
rect 31347 12804 31392 12832
rect 31386 12792 31392 12804
rect 31444 12792 31450 12844
rect 31938 12792 31944 12844
rect 31996 12832 32002 12844
rect 32769 12835 32827 12841
rect 32769 12832 32781 12835
rect 31996 12804 32781 12832
rect 31996 12792 32002 12804
rect 32769 12801 32781 12804
rect 32815 12801 32827 12835
rect 32769 12795 32827 12801
rect 24857 12767 24915 12773
rect 24857 12764 24869 12767
rect 24636 12736 24869 12764
rect 24636 12724 24642 12736
rect 24857 12733 24869 12736
rect 24903 12733 24915 12767
rect 24857 12727 24915 12733
rect 25041 12767 25099 12773
rect 25041 12733 25053 12767
rect 25087 12733 25099 12767
rect 25041 12727 25099 12733
rect 29917 12767 29975 12773
rect 29917 12733 29929 12767
rect 29963 12733 29975 12767
rect 29917 12727 29975 12733
rect 14182 12696 14188 12708
rect 10652 12668 14188 12696
rect 10652 12656 10658 12668
rect 14182 12656 14188 12668
rect 14240 12656 14246 12708
rect 29932 12696 29960 12727
rect 30006 12724 30012 12776
rect 30064 12764 30070 12776
rect 30101 12767 30159 12773
rect 30101 12764 30113 12767
rect 30064 12736 30113 12764
rect 30064 12724 30070 12736
rect 30101 12733 30113 12736
rect 30147 12733 30159 12767
rect 31202 12764 31208 12776
rect 31163 12736 31208 12764
rect 30101 12727 30159 12733
rect 31202 12724 31208 12736
rect 31260 12724 31266 12776
rect 31754 12696 31760 12708
rect 29932 12668 31760 12696
rect 31754 12656 31760 12668
rect 31812 12696 31818 12708
rect 32122 12696 32128 12708
rect 31812 12668 32128 12696
rect 31812 12656 31818 12668
rect 32122 12656 32128 12668
rect 32180 12656 32186 12708
rect 7006 12588 7012 12640
rect 7064 12628 7070 12640
rect 8297 12631 8355 12637
rect 8297 12628 8309 12631
rect 7064 12600 8309 12628
rect 7064 12588 7070 12600
rect 8297 12597 8309 12600
rect 8343 12597 8355 12631
rect 9122 12628 9128 12640
rect 9083 12600 9128 12628
rect 8297 12591 8355 12597
rect 9122 12588 9128 12600
rect 9180 12588 9186 12640
rect 11146 12588 11152 12640
rect 11204 12628 11210 12640
rect 11701 12631 11759 12637
rect 11701 12628 11713 12631
rect 11204 12600 11713 12628
rect 11204 12588 11210 12600
rect 11701 12597 11713 12600
rect 11747 12597 11759 12631
rect 11701 12591 11759 12597
rect 22189 12631 22247 12637
rect 22189 12597 22201 12631
rect 22235 12628 22247 12631
rect 22370 12628 22376 12640
rect 22235 12600 22376 12628
rect 22235 12597 22247 12600
rect 22189 12591 22247 12597
rect 22370 12588 22376 12600
rect 22428 12588 22434 12640
rect 24394 12628 24400 12640
rect 24355 12600 24400 12628
rect 24394 12588 24400 12600
rect 24452 12588 24458 12640
rect 1104 12538 37628 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 37628 12538
rect 1104 12464 37628 12486
rect 6365 12427 6423 12433
rect 6365 12393 6377 12427
rect 6411 12424 6423 12427
rect 6822 12424 6828 12436
rect 6411 12396 6828 12424
rect 6411 12393 6423 12396
rect 6365 12387 6423 12393
rect 6822 12384 6828 12396
rect 6880 12384 6886 12436
rect 8478 12384 8484 12436
rect 8536 12424 8542 12436
rect 8573 12427 8631 12433
rect 8573 12424 8585 12427
rect 8536 12396 8585 12424
rect 8536 12384 8542 12396
rect 8573 12393 8585 12396
rect 8619 12393 8631 12427
rect 13538 12424 13544 12436
rect 13499 12396 13544 12424
rect 8573 12387 8631 12393
rect 13538 12384 13544 12396
rect 13596 12384 13602 12436
rect 22833 12427 22891 12433
rect 22833 12393 22845 12427
rect 22879 12424 22891 12427
rect 22922 12424 22928 12436
rect 22879 12396 22928 12424
rect 22879 12393 22891 12396
rect 22833 12387 22891 12393
rect 22922 12384 22928 12396
rect 22980 12384 22986 12436
rect 26697 12427 26755 12433
rect 26697 12393 26709 12427
rect 26743 12424 26755 12427
rect 30190 12424 30196 12436
rect 26743 12396 30196 12424
rect 26743 12393 26755 12396
rect 26697 12387 26755 12393
rect 8294 12316 8300 12368
rect 8352 12356 8358 12368
rect 9398 12356 9404 12368
rect 8352 12328 9404 12356
rect 8352 12316 8358 12328
rect 9398 12316 9404 12328
rect 9456 12356 9462 12368
rect 11054 12356 11060 12368
rect 9456 12328 11060 12356
rect 9456 12316 9462 12328
rect 6546 12248 6552 12300
rect 6604 12288 6610 12300
rect 6825 12291 6883 12297
rect 6825 12288 6837 12291
rect 6604 12260 6837 12288
rect 6604 12248 6610 12260
rect 6825 12257 6837 12260
rect 6871 12257 6883 12291
rect 6825 12251 6883 12257
rect 8570 12248 8576 12300
rect 8628 12288 8634 12300
rect 9692 12297 9720 12328
rect 11054 12316 11060 12328
rect 11112 12316 11118 12368
rect 24578 12316 24584 12368
rect 24636 12356 24642 12368
rect 24636 12328 25084 12356
rect 24636 12316 24642 12328
rect 9677 12291 9735 12297
rect 8628 12260 9628 12288
rect 8628 12248 8634 12260
rect 9600 12232 9628 12260
rect 9677 12257 9689 12291
rect 9723 12257 9735 12291
rect 9677 12251 9735 12257
rect 11793 12291 11851 12297
rect 11793 12257 11805 12291
rect 11839 12288 11851 12291
rect 12434 12288 12440 12300
rect 11839 12260 12440 12288
rect 11839 12257 11851 12260
rect 11793 12251 11851 12257
rect 12434 12248 12440 12260
rect 12492 12248 12498 12300
rect 21085 12291 21143 12297
rect 21085 12257 21097 12291
rect 21131 12288 21143 12291
rect 22094 12288 22100 12300
rect 21131 12260 22100 12288
rect 21131 12257 21143 12260
rect 21085 12251 21143 12257
rect 22094 12248 22100 12260
rect 22152 12248 22158 12300
rect 23106 12248 23112 12300
rect 23164 12288 23170 12300
rect 23937 12291 23995 12297
rect 23937 12288 23949 12291
rect 23164 12260 23949 12288
rect 23164 12248 23170 12260
rect 23937 12257 23949 12260
rect 23983 12288 23995 12291
rect 24762 12288 24768 12300
rect 23983 12260 24768 12288
rect 23983 12257 23995 12260
rect 23937 12251 23995 12257
rect 24762 12248 24768 12260
rect 24820 12248 24826 12300
rect 24854 12248 24860 12300
rect 24912 12288 24918 12300
rect 24949 12291 25007 12297
rect 24949 12288 24961 12291
rect 24912 12260 24961 12288
rect 24912 12248 24918 12260
rect 24949 12257 24961 12260
rect 24995 12257 25007 12291
rect 25056 12288 25084 12328
rect 26712 12288 26740 12387
rect 30190 12384 30196 12396
rect 30248 12384 30254 12436
rect 31386 12384 31392 12436
rect 31444 12424 31450 12436
rect 31573 12427 31631 12433
rect 31573 12424 31585 12427
rect 31444 12396 31585 12424
rect 31444 12384 31450 12396
rect 31573 12393 31585 12396
rect 31619 12393 31631 12427
rect 31573 12387 31631 12393
rect 28902 12316 28908 12368
rect 28960 12356 28966 12368
rect 30650 12356 30656 12368
rect 28960 12328 30656 12356
rect 28960 12316 28966 12328
rect 30650 12316 30656 12328
rect 30708 12316 30714 12368
rect 34514 12356 34520 12368
rect 32048 12328 34520 12356
rect 25056 12260 26740 12288
rect 27157 12291 27215 12297
rect 24949 12251 25007 12257
rect 27157 12257 27169 12291
rect 27203 12288 27215 12291
rect 28074 12288 28080 12300
rect 27203 12260 28080 12288
rect 27203 12257 27215 12260
rect 27157 12251 27215 12257
rect 28074 12248 28080 12260
rect 28132 12248 28138 12300
rect 30668 12288 30696 12316
rect 32048 12300 32076 12328
rect 34514 12316 34520 12328
rect 34572 12316 34578 12368
rect 32030 12288 32036 12300
rect 30576 12260 30696 12288
rect 31991 12260 32036 12288
rect 6178 12220 6184 12232
rect 6139 12192 6184 12220
rect 6178 12180 6184 12192
rect 6236 12180 6242 12232
rect 9490 12220 9496 12232
rect 9451 12192 9496 12220
rect 9490 12180 9496 12192
rect 9548 12180 9554 12232
rect 9582 12180 9588 12232
rect 9640 12220 9646 12232
rect 10505 12223 10563 12229
rect 10505 12220 10517 12223
rect 9640 12192 10517 12220
rect 9640 12180 9646 12192
rect 10505 12189 10517 12192
rect 10551 12189 10563 12223
rect 11146 12220 11152 12232
rect 11107 12192 11152 12220
rect 10505 12183 10563 12189
rect 11146 12180 11152 12192
rect 11204 12180 11210 12232
rect 14458 12220 14464 12232
rect 14419 12192 14464 12220
rect 14458 12180 14464 12192
rect 14516 12180 14522 12232
rect 23661 12223 23719 12229
rect 23661 12189 23673 12223
rect 23707 12220 23719 12223
rect 24394 12220 24400 12232
rect 23707 12192 24400 12220
rect 23707 12189 23719 12192
rect 23661 12183 23719 12189
rect 24394 12180 24400 12192
rect 24452 12180 24458 12232
rect 28905 12223 28963 12229
rect 28905 12189 28917 12223
rect 28951 12220 28963 12223
rect 29822 12220 29828 12232
rect 28951 12192 29828 12220
rect 28951 12189 28963 12192
rect 28905 12183 28963 12189
rect 29822 12180 29828 12192
rect 29880 12180 29886 12232
rect 29914 12180 29920 12232
rect 29972 12220 29978 12232
rect 30576 12229 30604 12260
rect 32030 12248 32036 12260
rect 32088 12248 32094 12300
rect 32125 12291 32183 12297
rect 32125 12257 32137 12291
rect 32171 12288 32183 12291
rect 33321 12291 33379 12297
rect 33321 12288 33333 12291
rect 32171 12260 33333 12288
rect 32171 12257 32183 12260
rect 32125 12251 32183 12257
rect 33321 12257 33333 12260
rect 33367 12257 33379 12291
rect 33321 12251 33379 12257
rect 30561 12223 30619 12229
rect 29972 12192 30017 12220
rect 29972 12180 29978 12192
rect 30561 12189 30573 12223
rect 30607 12189 30619 12223
rect 30561 12183 30619 12189
rect 30926 12180 30932 12232
rect 30984 12220 30990 12232
rect 30984 12216 32076 12220
rect 32140 12216 32168 12251
rect 30984 12192 32168 12216
rect 30984 12180 30990 12192
rect 32048 12188 32168 12192
rect 32214 12180 32220 12232
rect 32272 12220 32278 12232
rect 34149 12223 34207 12229
rect 34149 12220 34161 12223
rect 32272 12192 34161 12220
rect 32272 12180 32278 12192
rect 34149 12189 34161 12192
rect 34195 12189 34207 12223
rect 34149 12183 34207 12189
rect 34790 12180 34796 12232
rect 34848 12220 34854 12232
rect 34885 12223 34943 12229
rect 34885 12220 34897 12223
rect 34848 12192 34897 12220
rect 34848 12180 34854 12192
rect 34885 12189 34897 12192
rect 34931 12189 34943 12223
rect 34885 12183 34943 12189
rect 7098 12152 7104 12164
rect 7059 12124 7104 12152
rect 7098 12112 7104 12124
rect 7156 12112 7162 12164
rect 7834 12112 7840 12164
rect 7892 12112 7898 12164
rect 12069 12155 12127 12161
rect 12069 12121 12081 12155
rect 12115 12121 12127 12155
rect 14369 12155 14427 12161
rect 14369 12152 14381 12155
rect 13294 12124 14381 12152
rect 12069 12115 12127 12121
rect 14369 12121 14381 12124
rect 14415 12121 14427 12155
rect 14369 12115 14427 12121
rect 21361 12155 21419 12161
rect 21361 12121 21373 12155
rect 21407 12152 21419 12155
rect 21450 12152 21456 12164
rect 21407 12124 21456 12152
rect 21407 12121 21419 12124
rect 21361 12115 21419 12121
rect 8662 12044 8668 12096
rect 8720 12084 8726 12096
rect 9125 12087 9183 12093
rect 9125 12084 9137 12087
rect 8720 12056 9137 12084
rect 8720 12044 8726 12056
rect 9125 12053 9137 12056
rect 9171 12053 9183 12087
rect 9125 12047 9183 12053
rect 9585 12087 9643 12093
rect 9585 12053 9597 12087
rect 9631 12084 9643 12087
rect 9674 12084 9680 12096
rect 9631 12056 9680 12084
rect 9631 12053 9643 12056
rect 9585 12047 9643 12053
rect 9674 12044 9680 12056
rect 9732 12044 9738 12096
rect 10597 12087 10655 12093
rect 10597 12053 10609 12087
rect 10643 12084 10655 12087
rect 10870 12084 10876 12096
rect 10643 12056 10876 12084
rect 10643 12053 10655 12056
rect 10597 12047 10655 12053
rect 10870 12044 10876 12056
rect 10928 12044 10934 12096
rect 11333 12087 11391 12093
rect 11333 12053 11345 12087
rect 11379 12084 11391 12087
rect 12084 12084 12112 12115
rect 21450 12112 21456 12124
rect 21508 12112 21514 12164
rect 22370 12112 22376 12164
rect 22428 12112 22434 12164
rect 24026 12112 24032 12164
rect 24084 12152 24090 12164
rect 25225 12155 25283 12161
rect 25225 12152 25237 12155
rect 24084 12124 25237 12152
rect 24084 12112 24090 12124
rect 25225 12121 25237 12124
rect 25271 12121 25283 12155
rect 27338 12152 27344 12164
rect 26450 12124 27344 12152
rect 25225 12115 25283 12121
rect 27338 12112 27344 12124
rect 27396 12112 27402 12164
rect 28198 12124 28580 12152
rect 23290 12084 23296 12096
rect 11379 12056 12112 12084
rect 23251 12056 23296 12084
rect 11379 12053 11391 12056
rect 11333 12047 11391 12053
rect 23290 12044 23296 12056
rect 23348 12044 23354 12096
rect 23750 12084 23756 12096
rect 23711 12056 23756 12084
rect 23750 12044 23756 12056
rect 23808 12044 23814 12096
rect 28552 12084 28580 12124
rect 28626 12112 28632 12164
rect 28684 12152 28690 12164
rect 30469 12155 30527 12161
rect 30469 12152 30481 12155
rect 28684 12124 28729 12152
rect 28828 12124 30481 12152
rect 28684 12112 28690 12124
rect 28828 12084 28856 12124
rect 30469 12121 30481 12124
rect 30515 12121 30527 12155
rect 33134 12152 33140 12164
rect 33095 12124 33140 12152
rect 30469 12115 30527 12121
rect 33134 12112 33140 12124
rect 33192 12112 33198 12164
rect 28552 12056 28856 12084
rect 29546 12044 29552 12096
rect 29604 12084 29610 12096
rect 29733 12087 29791 12093
rect 29733 12084 29745 12087
rect 29604 12056 29745 12084
rect 29604 12044 29610 12056
rect 29733 12053 29745 12056
rect 29779 12053 29791 12087
rect 29733 12047 29791 12053
rect 30006 12044 30012 12096
rect 30064 12084 30070 12096
rect 31941 12087 31999 12093
rect 31941 12084 31953 12087
rect 30064 12056 31953 12084
rect 30064 12044 30070 12056
rect 31941 12053 31953 12056
rect 31987 12053 31999 12087
rect 32766 12084 32772 12096
rect 32727 12056 32772 12084
rect 31941 12047 31999 12053
rect 32766 12044 32772 12056
rect 32824 12044 32830 12096
rect 33226 12044 33232 12096
rect 33284 12084 33290 12096
rect 33962 12084 33968 12096
rect 33284 12056 33329 12084
rect 33923 12056 33968 12084
rect 33284 12044 33290 12056
rect 33962 12044 33968 12056
rect 34020 12044 34026 12096
rect 34974 12084 34980 12096
rect 34935 12056 34980 12084
rect 34974 12044 34980 12056
rect 35032 12044 35038 12096
rect 1104 11994 37628 12016
rect 1104 11942 4874 11994
rect 4926 11942 4938 11994
rect 4990 11942 5002 11994
rect 5054 11942 5066 11994
rect 5118 11942 5130 11994
rect 5182 11942 35594 11994
rect 35646 11942 35658 11994
rect 35710 11942 35722 11994
rect 35774 11942 35786 11994
rect 35838 11942 35850 11994
rect 35902 11942 37628 11994
rect 1104 11920 37628 11942
rect 6178 11840 6184 11892
rect 6236 11880 6242 11892
rect 6549 11883 6607 11889
rect 6549 11880 6561 11883
rect 6236 11852 6561 11880
rect 6236 11840 6242 11852
rect 6549 11849 6561 11852
rect 6595 11849 6607 11883
rect 7834 11880 7840 11892
rect 7795 11852 7840 11880
rect 6549 11843 6607 11849
rect 7834 11840 7840 11852
rect 7892 11840 7898 11892
rect 9122 11840 9128 11892
rect 9180 11880 9186 11892
rect 9401 11883 9459 11889
rect 9401 11880 9413 11883
rect 9180 11852 9413 11880
rect 9180 11840 9186 11852
rect 9401 11849 9413 11852
rect 9447 11849 9459 11883
rect 9401 11843 9459 11849
rect 9493 11883 9551 11889
rect 9493 11849 9505 11883
rect 9539 11880 9551 11883
rect 9674 11880 9680 11892
rect 9539 11852 9680 11880
rect 9539 11849 9551 11852
rect 9493 11843 9551 11849
rect 9674 11840 9680 11852
rect 9732 11880 9738 11892
rect 10226 11880 10232 11892
rect 9732 11852 10232 11880
rect 9732 11840 9738 11852
rect 10226 11840 10232 11852
rect 10284 11840 10290 11892
rect 10689 11883 10747 11889
rect 10689 11849 10701 11883
rect 10735 11880 10747 11883
rect 11238 11880 11244 11892
rect 10735 11852 11244 11880
rect 10735 11849 10747 11852
rect 10689 11843 10747 11849
rect 11238 11840 11244 11852
rect 11296 11880 11302 11892
rect 11882 11880 11888 11892
rect 11296 11852 11888 11880
rect 11296 11840 11302 11852
rect 11882 11840 11888 11852
rect 11940 11840 11946 11892
rect 24578 11880 24584 11892
rect 24539 11852 24584 11880
rect 24578 11840 24584 11852
rect 24636 11840 24642 11892
rect 27338 11840 27344 11892
rect 27396 11880 27402 11892
rect 28445 11883 28503 11889
rect 28445 11880 28457 11883
rect 27396 11852 28457 11880
rect 27396 11840 27402 11852
rect 28445 11849 28457 11852
rect 28491 11849 28503 11883
rect 29086 11880 29092 11892
rect 29047 11852 29092 11880
rect 28445 11843 28503 11849
rect 29086 11840 29092 11852
rect 29144 11840 29150 11892
rect 30006 11880 30012 11892
rect 29967 11852 30012 11880
rect 30006 11840 30012 11852
rect 30064 11840 30070 11892
rect 31389 11883 31447 11889
rect 31389 11849 31401 11883
rect 31435 11880 31447 11883
rect 32766 11880 32772 11892
rect 31435 11852 32772 11880
rect 31435 11849 31447 11852
rect 31389 11843 31447 11849
rect 32766 11840 32772 11852
rect 32824 11840 32830 11892
rect 33226 11840 33232 11892
rect 33284 11880 33290 11892
rect 34793 11883 34851 11889
rect 34793 11880 34805 11883
rect 33284 11852 34805 11880
rect 33284 11840 33290 11852
rect 34793 11849 34805 11852
rect 34839 11880 34851 11883
rect 36630 11880 36636 11892
rect 34839 11852 36636 11880
rect 34839 11849 34851 11852
rect 34793 11843 34851 11849
rect 36630 11840 36636 11852
rect 36688 11840 36694 11892
rect 9582 11772 9588 11824
rect 9640 11812 9646 11824
rect 13630 11812 13636 11824
rect 9640 11784 13636 11812
rect 9640 11772 9646 11784
rect 13630 11772 13636 11784
rect 13688 11812 13694 11824
rect 13725 11815 13783 11821
rect 13725 11812 13737 11815
rect 13688 11784 13737 11812
rect 13688 11772 13694 11784
rect 13725 11781 13737 11784
rect 13771 11781 13783 11815
rect 22186 11812 22192 11824
rect 13725 11775 13783 11781
rect 22020 11784 22192 11812
rect 6914 11704 6920 11756
rect 6972 11744 6978 11756
rect 6972 11716 7017 11744
rect 6972 11704 6978 11716
rect 7282 11704 7288 11756
rect 7340 11744 7346 11756
rect 7745 11747 7803 11753
rect 7745 11744 7757 11747
rect 7340 11716 7757 11744
rect 7340 11704 7346 11716
rect 7745 11713 7757 11716
rect 7791 11744 7803 11747
rect 7926 11744 7932 11756
rect 7791 11716 7932 11744
rect 7791 11713 7803 11716
rect 7745 11707 7803 11713
rect 7926 11704 7932 11716
rect 7984 11704 7990 11756
rect 8389 11747 8447 11753
rect 8389 11713 8401 11747
rect 8435 11744 8447 11747
rect 10781 11747 10839 11753
rect 8435 11716 9076 11744
rect 8435 11713 8447 11716
rect 8389 11707 8447 11713
rect 7006 11676 7012 11688
rect 6967 11648 7012 11676
rect 7006 11636 7012 11648
rect 7064 11636 7070 11688
rect 7190 11676 7196 11688
rect 7151 11648 7196 11676
rect 7190 11636 7196 11648
rect 7248 11636 7254 11688
rect 9048 11617 9076 11716
rect 10781 11713 10793 11747
rect 10827 11744 10839 11747
rect 12342 11744 12348 11756
rect 10827 11716 12348 11744
rect 10827 11713 10839 11716
rect 10781 11707 10839 11713
rect 12342 11704 12348 11716
rect 12400 11704 12406 11756
rect 12618 11744 12624 11756
rect 12579 11716 12624 11744
rect 12618 11704 12624 11716
rect 12676 11704 12682 11756
rect 13449 11747 13507 11753
rect 13449 11713 13461 11747
rect 13495 11744 13507 11747
rect 14734 11744 14740 11756
rect 13495 11716 14740 11744
rect 13495 11713 13507 11716
rect 13449 11707 13507 11713
rect 14734 11704 14740 11716
rect 14792 11744 14798 11756
rect 17862 11744 17868 11756
rect 14792 11716 17868 11744
rect 14792 11704 14798 11716
rect 17862 11704 17868 11716
rect 17920 11704 17926 11756
rect 22020 11753 22048 11784
rect 22186 11772 22192 11784
rect 22244 11772 22250 11824
rect 23014 11772 23020 11824
rect 23072 11772 23078 11824
rect 24762 11772 24768 11824
rect 24820 11812 24826 11824
rect 24820 11784 26004 11812
rect 24820 11772 24826 11784
rect 22005 11747 22063 11753
rect 22005 11713 22017 11747
rect 22051 11713 22063 11747
rect 22005 11707 22063 11713
rect 25314 11704 25320 11756
rect 25372 11744 25378 11756
rect 25777 11747 25835 11753
rect 25777 11744 25789 11747
rect 25372 11716 25789 11744
rect 25372 11704 25378 11716
rect 25777 11713 25789 11716
rect 25823 11713 25835 11747
rect 25777 11707 25835 11713
rect 9677 11679 9735 11685
rect 9677 11645 9689 11679
rect 9723 11676 9735 11679
rect 10594 11676 10600 11688
rect 9723 11648 10600 11676
rect 9723 11645 9735 11648
rect 9677 11639 9735 11645
rect 10594 11636 10600 11648
rect 10652 11636 10658 11688
rect 11790 11676 11796 11688
rect 11751 11648 11796 11676
rect 11790 11636 11796 11648
rect 11848 11636 11854 11688
rect 22278 11676 22284 11688
rect 22239 11648 22284 11676
rect 22278 11636 22284 11648
rect 22336 11636 22342 11688
rect 23750 11676 23756 11688
rect 23663 11648 23756 11676
rect 23750 11636 23756 11648
rect 23808 11676 23814 11688
rect 24670 11676 24676 11688
rect 23808 11648 24676 11676
rect 23808 11636 23814 11648
rect 24670 11636 24676 11648
rect 24728 11636 24734 11688
rect 24765 11679 24823 11685
rect 24765 11645 24777 11679
rect 24811 11645 24823 11679
rect 24765 11639 24823 11645
rect 9033 11611 9091 11617
rect 9033 11577 9045 11611
rect 9079 11577 9091 11611
rect 24780 11608 24808 11639
rect 25590 11636 25596 11688
rect 25648 11676 25654 11688
rect 25976 11685 26004 11784
rect 26602 11772 26608 11824
rect 26660 11812 26666 11824
rect 27522 11812 27528 11824
rect 26660 11784 27528 11812
rect 26660 11772 26666 11784
rect 27522 11772 27528 11784
rect 27580 11772 27586 11824
rect 31297 11815 31355 11821
rect 31297 11781 31309 11815
rect 31343 11812 31355 11815
rect 33594 11812 33600 11824
rect 31343 11784 33600 11812
rect 31343 11781 31355 11784
rect 31297 11775 31355 11781
rect 33594 11772 33600 11784
rect 33652 11772 33658 11824
rect 34974 11812 34980 11824
rect 34546 11784 34980 11812
rect 34974 11772 34980 11784
rect 35032 11772 35038 11824
rect 26142 11704 26148 11756
rect 26200 11744 26206 11756
rect 27433 11747 27491 11753
rect 27433 11744 27445 11747
rect 26200 11716 27445 11744
rect 26200 11704 26206 11716
rect 27433 11713 27445 11716
rect 27479 11713 27491 11747
rect 27433 11707 27491 11713
rect 27614 11704 27620 11756
rect 27672 11744 27678 11756
rect 28537 11747 28595 11753
rect 28537 11744 28549 11747
rect 27672 11716 28549 11744
rect 27672 11704 27678 11716
rect 28537 11713 28549 11716
rect 28583 11744 28595 11747
rect 28902 11744 28908 11756
rect 28583 11716 28908 11744
rect 28583 11713 28595 11716
rect 28537 11707 28595 11713
rect 28902 11704 28908 11716
rect 28960 11744 28966 11756
rect 29181 11747 29239 11753
rect 29181 11744 29193 11747
rect 28960 11716 29193 11744
rect 28960 11704 28966 11716
rect 29181 11713 29193 11716
rect 29227 11713 29239 11747
rect 30098 11744 30104 11756
rect 30059 11716 30104 11744
rect 29181 11707 29239 11713
rect 30098 11704 30104 11716
rect 30156 11704 30162 11756
rect 30742 11704 30748 11756
rect 30800 11744 30806 11756
rect 32493 11747 32551 11753
rect 32493 11744 32505 11747
rect 30800 11716 32505 11744
rect 30800 11704 30806 11716
rect 32493 11713 32505 11716
rect 32539 11713 32551 11747
rect 32493 11707 32551 11713
rect 25869 11679 25927 11685
rect 25869 11676 25881 11679
rect 25648 11648 25881 11676
rect 25648 11636 25654 11648
rect 25869 11645 25881 11648
rect 25915 11645 25927 11679
rect 25869 11639 25927 11645
rect 25961 11679 26019 11685
rect 25961 11645 25973 11679
rect 26007 11645 26019 11679
rect 26234 11676 26240 11688
rect 25961 11639 26019 11645
rect 26206 11636 26240 11676
rect 26292 11676 26298 11688
rect 27338 11676 27344 11688
rect 26292 11648 27344 11676
rect 26292 11636 26298 11648
rect 27338 11636 27344 11648
rect 27396 11636 27402 11688
rect 29917 11679 29975 11685
rect 29917 11645 29929 11679
rect 29963 11676 29975 11679
rect 30190 11676 30196 11688
rect 29963 11648 30196 11676
rect 29963 11645 29975 11648
rect 29917 11639 29975 11645
rect 30190 11636 30196 11648
rect 30248 11636 30254 11688
rect 31202 11676 31208 11688
rect 31115 11648 31208 11676
rect 31202 11636 31208 11648
rect 31260 11676 31266 11688
rect 32030 11676 32036 11688
rect 31260 11648 32036 11676
rect 31260 11636 31266 11648
rect 32030 11636 32036 11648
rect 32088 11636 32094 11688
rect 33042 11676 33048 11688
rect 33003 11648 33048 11676
rect 33042 11636 33048 11648
rect 33100 11636 33106 11688
rect 33318 11676 33324 11688
rect 33279 11648 33324 11676
rect 33318 11636 33324 11648
rect 33376 11636 33382 11688
rect 26206 11608 26234 11636
rect 24780 11580 26234 11608
rect 27893 11611 27951 11617
rect 9033 11571 9091 11577
rect 27893 11577 27905 11611
rect 27939 11608 27951 11611
rect 28994 11608 29000 11620
rect 27939 11580 29000 11608
rect 27939 11577 27951 11580
rect 27893 11571 27951 11577
rect 28994 11568 29000 11580
rect 29052 11568 29058 11620
rect 30469 11611 30527 11617
rect 30469 11577 30481 11611
rect 30515 11608 30527 11611
rect 32214 11608 32220 11620
rect 30515 11580 32220 11608
rect 30515 11577 30527 11580
rect 30469 11571 30527 11577
rect 32214 11568 32220 11580
rect 32272 11568 32278 11620
rect 8573 11543 8631 11549
rect 8573 11509 8585 11543
rect 8619 11540 8631 11543
rect 8754 11540 8760 11552
rect 8619 11512 8760 11540
rect 8619 11509 8631 11512
rect 8573 11503 8631 11509
rect 8754 11500 8760 11512
rect 8812 11500 8818 11552
rect 11146 11540 11152 11552
rect 11107 11512 11152 11540
rect 11146 11500 11152 11512
rect 11204 11500 11210 11552
rect 23842 11500 23848 11552
rect 23900 11540 23906 11552
rect 24213 11543 24271 11549
rect 24213 11540 24225 11543
rect 23900 11512 24225 11540
rect 23900 11500 23906 11512
rect 24213 11509 24225 11512
rect 24259 11509 24271 11543
rect 24213 11503 24271 11509
rect 24302 11500 24308 11552
rect 24360 11540 24366 11552
rect 25409 11543 25467 11549
rect 25409 11540 25421 11543
rect 24360 11512 25421 11540
rect 24360 11500 24366 11512
rect 25409 11509 25421 11512
rect 25455 11509 25467 11543
rect 31754 11540 31760 11552
rect 31715 11512 31760 11540
rect 25409 11503 25467 11509
rect 31754 11500 31760 11512
rect 31812 11500 31818 11552
rect 32398 11540 32404 11552
rect 32359 11512 32404 11540
rect 32398 11500 32404 11512
rect 32456 11500 32462 11552
rect 1104 11450 37628 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 37628 11450
rect 1104 11376 37628 11398
rect 7098 11296 7104 11348
rect 7156 11336 7162 11348
rect 7653 11339 7711 11345
rect 7653 11336 7665 11339
rect 7156 11308 7665 11336
rect 7156 11296 7162 11308
rect 7653 11305 7665 11308
rect 7699 11305 7711 11339
rect 11882 11336 11888 11348
rect 11843 11308 11888 11336
rect 7653 11299 7711 11305
rect 11882 11296 11888 11308
rect 11940 11296 11946 11348
rect 12342 11336 12348 11348
rect 12303 11308 12348 11336
rect 12342 11296 12348 11308
rect 12400 11296 12406 11348
rect 22278 11336 22284 11348
rect 22239 11308 22284 11336
rect 22278 11296 22284 11308
rect 22336 11296 22342 11348
rect 23014 11336 23020 11348
rect 22975 11308 23020 11336
rect 23014 11296 23020 11308
rect 23072 11296 23078 11348
rect 24026 11336 24032 11348
rect 23987 11308 24032 11336
rect 24026 11296 24032 11308
rect 24084 11296 24090 11348
rect 25314 11336 25320 11348
rect 25275 11308 25320 11336
rect 25314 11296 25320 11308
rect 25372 11296 25378 11348
rect 29825 11339 29883 11345
rect 29825 11305 29837 11339
rect 29871 11336 29883 11339
rect 30006 11336 30012 11348
rect 29871 11308 30012 11336
rect 29871 11305 29883 11308
rect 29825 11299 29883 11305
rect 30006 11296 30012 11308
rect 30064 11296 30070 11348
rect 31315 11339 31373 11345
rect 31315 11305 31327 11339
rect 31361 11336 31373 11339
rect 33962 11336 33968 11348
rect 31361 11308 33968 11336
rect 31361 11305 31373 11308
rect 31315 11299 31373 11305
rect 33962 11296 33968 11308
rect 34020 11296 34026 11348
rect 24946 11268 24952 11280
rect 12636 11240 12940 11268
rect 9766 11160 9772 11212
rect 9824 11200 9830 11212
rect 12636 11200 12664 11240
rect 12802 11200 12808 11212
rect 9824 11172 12664 11200
rect 12763 11172 12808 11200
rect 9824 11160 9830 11172
rect 12802 11160 12808 11172
rect 12860 11160 12866 11212
rect 12912 11209 12940 11240
rect 24780 11240 24952 11268
rect 12897 11203 12955 11209
rect 12897 11169 12909 11203
rect 12943 11169 12955 11203
rect 23290 11200 23296 11212
rect 12897 11163 12955 11169
rect 22480 11172 23296 11200
rect 6549 11135 6607 11141
rect 6549 11101 6561 11135
rect 6595 11132 6607 11135
rect 6638 11132 6644 11144
rect 6595 11104 6644 11132
rect 6595 11101 6607 11104
rect 6549 11095 6607 11101
rect 6638 11092 6644 11104
rect 6696 11092 6702 11144
rect 7837 11135 7895 11141
rect 7837 11101 7849 11135
rect 7883 11132 7895 11135
rect 8662 11132 8668 11144
rect 7883 11104 8668 11132
rect 7883 11101 7895 11104
rect 7837 11095 7895 11101
rect 8662 11092 8668 11104
rect 8720 11092 8726 11144
rect 9493 11135 9551 11141
rect 9493 11101 9505 11135
rect 9539 11132 9551 11135
rect 9582 11132 9588 11144
rect 9539 11104 9588 11132
rect 9539 11101 9551 11104
rect 9493 11095 9551 11101
rect 9582 11092 9588 11104
rect 9640 11092 9646 11144
rect 10134 11132 10140 11144
rect 10095 11104 10140 11132
rect 10134 11092 10140 11104
rect 10192 11092 10198 11144
rect 13725 11135 13783 11141
rect 13725 11101 13737 11135
rect 13771 11132 13783 11135
rect 14458 11132 14464 11144
rect 13771 11104 14464 11132
rect 13771 11101 13783 11104
rect 13725 11095 13783 11101
rect 14458 11092 14464 11104
rect 14516 11132 14522 11144
rect 17218 11132 17224 11144
rect 14516 11104 17224 11132
rect 14516 11092 14522 11104
rect 17218 11092 17224 11104
rect 17276 11092 17282 11144
rect 22480 11141 22508 11172
rect 23290 11160 23296 11172
rect 23348 11160 23354 11212
rect 24578 11160 24584 11212
rect 24636 11200 24642 11212
rect 24780 11209 24808 11240
rect 24946 11228 24952 11240
rect 25004 11268 25010 11280
rect 25004 11240 26924 11268
rect 25004 11228 25010 11240
rect 24765 11203 24823 11209
rect 24765 11200 24777 11203
rect 24636 11172 24777 11200
rect 24636 11160 24642 11172
rect 24765 11169 24777 11172
rect 24811 11169 24823 11203
rect 24765 11163 24823 11169
rect 24857 11203 24915 11209
rect 24857 11169 24869 11203
rect 24903 11200 24915 11203
rect 26602 11200 26608 11212
rect 24903 11172 26608 11200
rect 24903 11169 24915 11172
rect 24857 11163 24915 11169
rect 26602 11160 26608 11172
rect 26660 11160 26666 11212
rect 26896 11209 26924 11240
rect 27338 11228 27344 11280
rect 27396 11268 27402 11280
rect 30190 11268 30196 11280
rect 27396 11240 30196 11268
rect 27396 11228 27402 11240
rect 27632 11209 27660 11240
rect 30190 11228 30196 11240
rect 30248 11228 30254 11280
rect 33594 11228 33600 11280
rect 33652 11268 33658 11280
rect 33781 11271 33839 11277
rect 33781 11268 33793 11271
rect 33652 11240 33793 11268
rect 33652 11228 33658 11240
rect 33781 11237 33793 11240
rect 33827 11237 33839 11271
rect 33781 11231 33839 11237
rect 26881 11203 26939 11209
rect 26881 11169 26893 11203
rect 26927 11169 26939 11203
rect 26881 11163 26939 11169
rect 27617 11203 27675 11209
rect 27617 11169 27629 11203
rect 27663 11169 27675 11203
rect 27617 11163 27675 11169
rect 22465 11135 22523 11141
rect 22465 11101 22477 11135
rect 22511 11101 22523 11135
rect 22465 11095 22523 11101
rect 22830 11092 22836 11144
rect 22888 11132 22894 11144
rect 22925 11135 22983 11141
rect 22925 11132 22937 11135
rect 22888 11104 22937 11132
rect 22888 11092 22894 11104
rect 22925 11101 22937 11104
rect 22971 11101 22983 11135
rect 23842 11132 23848 11144
rect 23803 11104 23848 11132
rect 22925 11095 22983 11101
rect 23842 11092 23848 11104
rect 23900 11092 23906 11144
rect 26896 11132 26924 11163
rect 29822 11160 29828 11212
rect 29880 11200 29886 11212
rect 31573 11203 31631 11209
rect 31573 11200 31585 11203
rect 29880 11172 31585 11200
rect 29880 11160 29886 11172
rect 31573 11169 31585 11172
rect 31619 11200 31631 11203
rect 32033 11203 32091 11209
rect 32033 11200 32045 11203
rect 31619 11172 32045 11200
rect 31619 11169 31631 11172
rect 31573 11163 31631 11169
rect 32033 11169 32045 11172
rect 32079 11200 32091 11203
rect 33042 11200 33048 11212
rect 32079 11172 33048 11200
rect 32079 11169 32091 11172
rect 32033 11163 32091 11169
rect 33042 11160 33048 11172
rect 33100 11160 33106 11212
rect 26896 11104 28764 11132
rect 10410 11064 10416 11076
rect 10371 11036 10416 11064
rect 10410 11024 10416 11036
rect 10468 11024 10474 11076
rect 10870 11024 10876 11076
rect 10928 11024 10934 11076
rect 13538 11024 13544 11076
rect 13596 11064 13602 11076
rect 13633 11067 13691 11073
rect 13633 11064 13645 11067
rect 13596 11036 13645 11064
rect 13596 11024 13602 11036
rect 13633 11033 13645 11036
rect 13679 11033 13691 11067
rect 13633 11027 13691 11033
rect 24670 11024 24676 11076
rect 24728 11064 24734 11076
rect 24949 11067 25007 11073
rect 24949 11064 24961 11067
rect 24728 11036 24961 11064
rect 24728 11024 24734 11036
rect 24949 11033 24961 11036
rect 24995 11033 25007 11067
rect 24949 11027 25007 11033
rect 25590 11024 25596 11076
rect 25648 11064 25654 11076
rect 26142 11064 26148 11076
rect 25648 11036 26148 11064
rect 25648 11024 25654 11036
rect 26142 11024 26148 11036
rect 26200 11064 26206 11076
rect 26605 11067 26663 11073
rect 26605 11064 26617 11067
rect 26200 11036 26617 11064
rect 26200 11024 26206 11036
rect 26605 11033 26617 11036
rect 26651 11033 26663 11067
rect 26605 11027 26663 11033
rect 26697 11067 26755 11073
rect 26697 11033 26709 11067
rect 26743 11064 26755 11067
rect 27706 11064 27712 11076
rect 26743 11036 27568 11064
rect 27667 11036 27712 11064
rect 26743 11033 26755 11036
rect 26697 11027 26755 11033
rect 6362 10996 6368 11008
rect 6323 10968 6368 10996
rect 6362 10956 6368 10968
rect 6420 10956 6426 11008
rect 9490 10956 9496 11008
rect 9548 10996 9554 11008
rect 9585 10999 9643 11005
rect 9585 10996 9597 10999
rect 9548 10968 9597 10996
rect 9548 10956 9554 10968
rect 9585 10965 9597 10968
rect 9631 10965 9643 10999
rect 12710 10996 12716 11008
rect 12671 10968 12716 10996
rect 9585 10959 9643 10965
rect 12710 10956 12716 10968
rect 12768 10956 12774 11008
rect 26234 10956 26240 11008
rect 26292 10996 26298 11008
rect 27540 10996 27568 11036
rect 27706 11024 27712 11036
rect 27764 11024 27770 11076
rect 27801 11067 27859 11073
rect 27801 11033 27813 11067
rect 27847 11064 27859 11067
rect 28074 11064 28080 11076
rect 27847 11036 28080 11064
rect 27847 11033 27859 11036
rect 27801 11027 27859 11033
rect 27816 10996 27844 11027
rect 28074 11024 28080 11036
rect 28132 11024 28138 11076
rect 28736 11073 28764 11104
rect 34330 11092 34336 11144
rect 34388 11132 34394 11144
rect 35069 11135 35127 11141
rect 35069 11132 35081 11135
rect 34388 11104 35081 11132
rect 34388 11092 34394 11104
rect 35069 11101 35081 11104
rect 35115 11101 35127 11135
rect 35069 11095 35127 11101
rect 28721 11067 28779 11073
rect 28721 11033 28733 11067
rect 28767 11064 28779 11067
rect 28902 11064 28908 11076
rect 28767 11036 28908 11064
rect 28767 11033 28779 11036
rect 28721 11027 28779 11033
rect 28902 11024 28908 11036
rect 28960 11024 28966 11076
rect 29089 11067 29147 11073
rect 29089 11033 29101 11067
rect 29135 11064 29147 11067
rect 32306 11064 32312 11076
rect 29135 11036 30052 11064
rect 30866 11036 31248 11064
rect 29135 11033 29147 11036
rect 29089 11027 29147 11033
rect 28166 10996 28172 11008
rect 26292 10968 26337 10996
rect 27540 10968 27844 10996
rect 28127 10968 28172 10996
rect 26292 10956 26298 10968
rect 28166 10956 28172 10968
rect 28224 10956 28230 11008
rect 30024 10996 30052 11036
rect 30926 10996 30932 11008
rect 30024 10968 30932 10996
rect 30926 10956 30932 10968
rect 30984 10956 30990 11008
rect 31220 10996 31248 11036
rect 31404 11036 32168 11064
rect 32267 11036 32312 11064
rect 31404 10996 31432 11036
rect 31220 10968 31432 10996
rect 32140 10996 32168 11036
rect 32306 11024 32312 11036
rect 32364 11024 32370 11076
rect 34977 11067 35035 11073
rect 34977 11064 34989 11067
rect 33534 11036 34989 11064
rect 34977 11033 34989 11036
rect 35023 11033 35035 11067
rect 34977 11027 35035 11033
rect 33686 10996 33692 11008
rect 32140 10968 33692 10996
rect 33686 10956 33692 10968
rect 33744 10956 33750 11008
rect 1104 10906 37628 10928
rect 1104 10854 4874 10906
rect 4926 10854 4938 10906
rect 4990 10854 5002 10906
rect 5054 10854 5066 10906
rect 5118 10854 5130 10906
rect 5182 10854 35594 10906
rect 35646 10854 35658 10906
rect 35710 10854 35722 10906
rect 35774 10854 35786 10906
rect 35838 10854 35850 10906
rect 35902 10854 37628 10906
rect 1104 10832 37628 10854
rect 1854 10752 1860 10804
rect 1912 10792 1918 10804
rect 8386 10792 8392 10804
rect 1912 10764 8392 10792
rect 1912 10752 1918 10764
rect 8386 10752 8392 10764
rect 8444 10752 8450 10804
rect 10134 10792 10140 10804
rect 8496 10764 10140 10792
rect 6546 10684 6552 10736
rect 6604 10724 6610 10736
rect 8496 10724 8524 10764
rect 10134 10752 10140 10764
rect 10192 10752 10198 10804
rect 10226 10752 10232 10804
rect 10284 10792 10290 10804
rect 10284 10764 10329 10792
rect 10284 10752 10290 10764
rect 10410 10752 10416 10804
rect 10468 10792 10474 10804
rect 10689 10795 10747 10801
rect 10689 10792 10701 10795
rect 10468 10764 10701 10792
rect 10468 10752 10474 10764
rect 10689 10761 10701 10764
rect 10735 10761 10747 10795
rect 10689 10755 10747 10761
rect 24673 10795 24731 10801
rect 24673 10761 24685 10795
rect 24719 10792 24731 10795
rect 24762 10792 24768 10804
rect 24719 10764 24768 10792
rect 24719 10761 24731 10764
rect 24673 10755 24731 10761
rect 24762 10752 24768 10764
rect 24820 10752 24826 10804
rect 25869 10795 25927 10801
rect 25869 10761 25881 10795
rect 25915 10792 25927 10795
rect 26234 10792 26240 10804
rect 25915 10764 26240 10792
rect 25915 10761 25927 10764
rect 25869 10755 25927 10761
rect 26234 10752 26240 10764
rect 26292 10752 26298 10804
rect 29380 10764 29684 10792
rect 8754 10724 8760 10736
rect 6604 10696 8524 10724
rect 8715 10696 8760 10724
rect 6604 10684 6610 10696
rect 6917 10659 6975 10665
rect 6917 10625 6929 10659
rect 6963 10656 6975 10659
rect 7834 10656 7840 10668
rect 6963 10628 7840 10656
rect 6963 10625 6975 10628
rect 6917 10619 6975 10625
rect 7834 10616 7840 10628
rect 7892 10616 7898 10668
rect 7926 10616 7932 10668
rect 7984 10656 7990 10668
rect 8496 10665 8524 10696
rect 8754 10684 8760 10696
rect 8812 10684 8818 10736
rect 9490 10684 9496 10736
rect 9548 10684 9554 10736
rect 10152 10724 10180 10752
rect 11790 10724 11796 10736
rect 10152 10696 11796 10724
rect 11790 10684 11796 10696
rect 11848 10724 11854 10736
rect 24302 10724 24308 10736
rect 11848 10696 12204 10724
rect 11848 10684 11854 10696
rect 8481 10659 8539 10665
rect 7984 10628 8029 10656
rect 7984 10616 7990 10628
rect 8481 10625 8493 10659
rect 8527 10625 8539 10659
rect 8481 10619 8539 10625
rect 10873 10659 10931 10665
rect 10873 10625 10885 10659
rect 10919 10656 10931 10659
rect 11146 10656 11152 10668
rect 10919 10628 11152 10656
rect 10919 10625 10931 10628
rect 10873 10619 10931 10625
rect 11146 10616 11152 10628
rect 11204 10616 11210 10668
rect 12176 10665 12204 10696
rect 22756 10696 24308 10724
rect 12161 10659 12219 10665
rect 12161 10625 12173 10659
rect 12207 10625 12219 10659
rect 12161 10619 12219 10625
rect 13538 10616 13544 10668
rect 13596 10616 13602 10668
rect 17862 10656 17868 10668
rect 17823 10628 17868 10656
rect 17862 10616 17868 10628
rect 17920 10616 17926 10668
rect 22756 10665 22784 10696
rect 24302 10684 24308 10696
rect 24360 10684 24366 10736
rect 26970 10684 26976 10736
rect 27028 10724 27034 10736
rect 27433 10727 27491 10733
rect 27433 10724 27445 10727
rect 27028 10696 27445 10724
rect 27028 10684 27034 10696
rect 27433 10693 27445 10696
rect 27479 10693 27491 10727
rect 29380 10724 29408 10764
rect 29546 10724 29552 10736
rect 29118 10696 29408 10724
rect 29507 10696 29552 10724
rect 27433 10687 27491 10693
rect 29546 10684 29552 10696
rect 29604 10684 29610 10736
rect 29656 10724 29684 10764
rect 30098 10752 30104 10804
rect 30156 10792 30162 10804
rect 30285 10795 30343 10801
rect 30285 10792 30297 10795
rect 30156 10764 30297 10792
rect 30156 10752 30162 10764
rect 30285 10761 30297 10764
rect 30331 10761 30343 10795
rect 30285 10755 30343 10761
rect 30466 10752 30472 10804
rect 30524 10792 30530 10804
rect 30745 10795 30803 10801
rect 30745 10792 30757 10795
rect 30524 10764 30757 10792
rect 30524 10752 30530 10764
rect 30745 10761 30757 10764
rect 30791 10761 30803 10795
rect 30745 10755 30803 10761
rect 32493 10795 32551 10801
rect 32493 10761 32505 10795
rect 32539 10792 32551 10795
rect 33318 10792 33324 10804
rect 32539 10764 33324 10792
rect 32539 10761 32551 10764
rect 32493 10755 32551 10761
rect 33318 10752 33324 10764
rect 33376 10752 33382 10804
rect 33413 10795 33471 10801
rect 33413 10761 33425 10795
rect 33459 10792 33471 10795
rect 33594 10792 33600 10804
rect 33459 10764 33600 10792
rect 33459 10761 33471 10764
rect 33413 10755 33471 10761
rect 32398 10724 32404 10736
rect 29656 10696 32404 10724
rect 32398 10684 32404 10696
rect 32456 10684 32462 10736
rect 33134 10684 33140 10736
rect 33192 10724 33198 10736
rect 33428 10724 33456 10755
rect 33594 10752 33600 10764
rect 33652 10752 33658 10804
rect 33686 10752 33692 10804
rect 33744 10792 33750 10804
rect 34241 10795 34299 10801
rect 34241 10792 34253 10795
rect 33744 10764 34253 10792
rect 33744 10752 33750 10764
rect 34241 10761 34253 10764
rect 34287 10761 34299 10795
rect 34241 10755 34299 10761
rect 33192 10696 33456 10724
rect 33192 10684 33198 10696
rect 22741 10659 22799 10665
rect 22741 10625 22753 10659
rect 22787 10625 22799 10659
rect 22741 10619 22799 10625
rect 23569 10659 23627 10665
rect 23569 10625 23581 10659
rect 23615 10656 23627 10659
rect 24578 10656 24584 10668
rect 23615 10628 24584 10656
rect 23615 10625 23627 10628
rect 23569 10619 23627 10625
rect 24578 10616 24584 10628
rect 24636 10616 24642 10668
rect 24949 10659 25007 10665
rect 24949 10625 24961 10659
rect 24995 10656 25007 10659
rect 26050 10656 26056 10668
rect 24995 10628 26056 10656
rect 24995 10625 25007 10628
rect 24949 10619 25007 10625
rect 26050 10616 26056 10628
rect 26108 10656 26114 10668
rect 27062 10656 27068 10668
rect 26108 10628 27068 10656
rect 26108 10616 26114 10628
rect 27062 10616 27068 10628
rect 27120 10656 27126 10668
rect 27157 10659 27215 10665
rect 27157 10656 27169 10659
rect 27120 10628 27169 10656
rect 27120 10616 27126 10628
rect 27157 10625 27169 10628
rect 27203 10625 27215 10659
rect 27157 10619 27215 10625
rect 29822 10616 29828 10668
rect 29880 10656 29886 10668
rect 30650 10656 30656 10668
rect 29880 10628 29925 10656
rect 30611 10628 30656 10656
rect 29880 10616 29886 10628
rect 30650 10616 30656 10628
rect 30708 10616 30714 10668
rect 31386 10616 31392 10668
rect 31444 10656 31450 10668
rect 31665 10659 31723 10665
rect 31665 10656 31677 10659
rect 31444 10628 31677 10656
rect 31444 10616 31450 10628
rect 31665 10625 31677 10628
rect 31711 10625 31723 10659
rect 31665 10619 31723 10625
rect 32309 10659 32367 10665
rect 32309 10625 32321 10659
rect 32355 10656 32367 10659
rect 32355 10628 32996 10656
rect 32355 10625 32367 10628
rect 32309 10619 32367 10625
rect 7006 10588 7012 10600
rect 6967 10560 7012 10588
rect 7006 10548 7012 10560
rect 7064 10548 7070 10600
rect 7193 10591 7251 10597
rect 7193 10557 7205 10591
rect 7239 10588 7251 10591
rect 8294 10588 8300 10600
rect 7239 10560 8300 10588
rect 7239 10557 7251 10560
rect 7193 10551 7251 10557
rect 8294 10548 8300 10560
rect 8352 10548 8358 10600
rect 11790 10548 11796 10600
rect 11848 10588 11854 10600
rect 12437 10591 12495 10597
rect 12437 10588 12449 10591
rect 11848 10560 12449 10588
rect 11848 10548 11854 10560
rect 12437 10557 12449 10560
rect 12483 10557 12495 10591
rect 12437 10551 12495 10557
rect 17681 10591 17739 10597
rect 17681 10557 17693 10591
rect 17727 10588 17739 10591
rect 18414 10588 18420 10600
rect 17727 10560 18420 10588
rect 17727 10557 17739 10560
rect 17681 10551 17739 10557
rect 18414 10548 18420 10560
rect 18472 10548 18478 10600
rect 25958 10588 25964 10600
rect 25919 10560 25964 10588
rect 25958 10548 25964 10560
rect 26016 10548 26022 10600
rect 26145 10591 26203 10597
rect 26145 10557 26157 10591
rect 26191 10588 26203 10591
rect 26234 10588 26240 10600
rect 26191 10560 26240 10588
rect 26191 10557 26203 10560
rect 26145 10551 26203 10557
rect 26234 10548 26240 10560
rect 26292 10588 26298 10600
rect 26970 10588 26976 10600
rect 26292 10560 26976 10588
rect 26292 10548 26298 10560
rect 26970 10548 26976 10560
rect 27028 10548 27034 10600
rect 28077 10591 28135 10597
rect 28077 10557 28089 10591
rect 28123 10588 28135 10591
rect 28810 10588 28816 10600
rect 28123 10560 28816 10588
rect 28123 10557 28135 10560
rect 28077 10551 28135 10557
rect 28810 10548 28816 10560
rect 28868 10588 28874 10600
rect 29454 10588 29460 10600
rect 28868 10560 29460 10588
rect 28868 10548 28874 10560
rect 29454 10548 29460 10560
rect 29512 10548 29518 10600
rect 30834 10588 30840 10600
rect 30795 10560 30840 10588
rect 30834 10548 30840 10560
rect 30892 10548 30898 10600
rect 6549 10523 6607 10529
rect 6549 10489 6561 10523
rect 6595 10520 6607 10523
rect 6638 10520 6644 10532
rect 6595 10492 6644 10520
rect 6595 10489 6607 10492
rect 6549 10483 6607 10489
rect 6638 10480 6644 10492
rect 6696 10480 6702 10532
rect 32968 10529 32996 10628
rect 33226 10616 33232 10668
rect 33284 10656 33290 10668
rect 33321 10659 33379 10665
rect 33321 10656 33333 10659
rect 33284 10628 33333 10656
rect 33284 10616 33290 10628
rect 33321 10625 33333 10628
rect 33367 10625 33379 10659
rect 33321 10619 33379 10625
rect 33686 10616 33692 10668
rect 33744 10656 33750 10668
rect 34330 10656 34336 10668
rect 33744 10628 34336 10656
rect 33744 10616 33750 10628
rect 34330 10616 34336 10628
rect 34388 10616 34394 10668
rect 33505 10591 33563 10597
rect 33505 10557 33517 10591
rect 33551 10557 33563 10591
rect 33505 10551 33563 10557
rect 32953 10523 33011 10529
rect 32953 10489 32965 10523
rect 32999 10489 33011 10523
rect 32953 10483 33011 10489
rect 7650 10412 7656 10464
rect 7708 10452 7714 10464
rect 7837 10455 7895 10461
rect 7837 10452 7849 10455
rect 7708 10424 7849 10452
rect 7708 10412 7714 10424
rect 7837 10421 7849 10424
rect 7883 10421 7895 10455
rect 13906 10452 13912 10464
rect 13867 10424 13912 10452
rect 7837 10415 7895 10421
rect 13906 10412 13912 10424
rect 13964 10412 13970 10464
rect 22554 10452 22560 10464
rect 22515 10424 22560 10452
rect 22554 10412 22560 10424
rect 22612 10412 22618 10464
rect 23106 10412 23112 10464
rect 23164 10452 23170 10464
rect 23293 10455 23351 10461
rect 23293 10452 23305 10455
rect 23164 10424 23305 10452
rect 23164 10412 23170 10424
rect 23293 10421 23305 10424
rect 23339 10421 23351 10455
rect 23293 10415 23351 10421
rect 24946 10412 24952 10464
rect 25004 10452 25010 10464
rect 25501 10455 25559 10461
rect 25501 10452 25513 10455
rect 25004 10424 25513 10452
rect 25004 10412 25010 10424
rect 25501 10421 25513 10424
rect 25547 10421 25559 10455
rect 25501 10415 25559 10421
rect 30374 10412 30380 10464
rect 30432 10452 30438 10464
rect 31481 10455 31539 10461
rect 31481 10452 31493 10455
rect 30432 10424 31493 10452
rect 30432 10412 30438 10424
rect 31481 10421 31493 10424
rect 31527 10421 31539 10455
rect 31481 10415 31539 10421
rect 31846 10412 31852 10464
rect 31904 10452 31910 10464
rect 32674 10452 32680 10464
rect 31904 10424 32680 10452
rect 31904 10412 31910 10424
rect 32674 10412 32680 10424
rect 32732 10452 32738 10464
rect 33520 10452 33548 10551
rect 32732 10424 33548 10452
rect 32732 10412 32738 10424
rect 1104 10362 37628 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 37628 10362
rect 1104 10288 37628 10310
rect 11790 10248 11796 10260
rect 11751 10220 11796 10248
rect 11790 10208 11796 10220
rect 11848 10208 11854 10260
rect 24029 10251 24087 10257
rect 24029 10217 24041 10251
rect 24075 10248 24087 10251
rect 25590 10248 25596 10260
rect 24075 10220 25596 10248
rect 24075 10217 24087 10220
rect 24029 10211 24087 10217
rect 25590 10208 25596 10220
rect 25648 10208 25654 10260
rect 28626 10208 28632 10260
rect 28684 10248 28690 10260
rect 28905 10251 28963 10257
rect 28905 10248 28917 10251
rect 28684 10220 28917 10248
rect 28684 10208 28690 10220
rect 28905 10217 28917 10220
rect 28951 10217 28963 10251
rect 28905 10211 28963 10217
rect 29733 10251 29791 10257
rect 29733 10217 29745 10251
rect 29779 10248 29791 10251
rect 29914 10248 29920 10260
rect 29779 10220 29920 10248
rect 29779 10217 29791 10220
rect 29733 10211 29791 10217
rect 29914 10208 29920 10220
rect 29972 10208 29978 10260
rect 30558 10208 30564 10260
rect 30616 10248 30622 10260
rect 31297 10251 31355 10257
rect 31297 10248 31309 10251
rect 30616 10220 31309 10248
rect 30616 10208 30622 10220
rect 31297 10217 31309 10220
rect 31343 10248 31355 10251
rect 31846 10248 31852 10260
rect 31343 10220 31852 10248
rect 31343 10217 31355 10220
rect 31297 10211 31355 10217
rect 31846 10208 31852 10220
rect 31904 10208 31910 10260
rect 32306 10208 32312 10260
rect 32364 10248 32370 10260
rect 33321 10251 33379 10257
rect 33321 10248 33333 10251
rect 32364 10220 33333 10248
rect 32364 10208 32370 10220
rect 33321 10217 33333 10220
rect 33367 10217 33379 10251
rect 33321 10211 33379 10217
rect 8386 10140 8392 10192
rect 8444 10180 8450 10192
rect 8444 10152 9260 10180
rect 8444 10140 8450 10152
rect 6089 10115 6147 10121
rect 6089 10081 6101 10115
rect 6135 10112 6147 10115
rect 6454 10112 6460 10124
rect 6135 10084 6460 10112
rect 6135 10081 6147 10084
rect 6089 10075 6147 10081
rect 6454 10072 6460 10084
rect 6512 10112 6518 10124
rect 9125 10115 9183 10121
rect 9125 10112 9137 10115
rect 6512 10084 9137 10112
rect 6512 10072 6518 10084
rect 9125 10081 9137 10084
rect 9171 10081 9183 10115
rect 9232 10112 9260 10152
rect 25958 10140 25964 10192
rect 26016 10180 26022 10192
rect 26329 10183 26387 10189
rect 26329 10180 26341 10183
rect 26016 10152 26341 10180
rect 26016 10140 26022 10152
rect 26329 10149 26341 10152
rect 26375 10180 26387 10183
rect 27706 10180 27712 10192
rect 26375 10152 27712 10180
rect 26375 10149 26387 10152
rect 26329 10143 26387 10149
rect 27706 10140 27712 10152
rect 27764 10140 27770 10192
rect 12710 10112 12716 10124
rect 9232 10084 12388 10112
rect 12671 10084 12716 10112
rect 9125 10075 9183 10081
rect 8386 10044 8392 10056
rect 8347 10016 8392 10044
rect 8386 10004 8392 10016
rect 8444 10004 8450 10056
rect 11609 10047 11667 10053
rect 11609 10013 11621 10047
rect 11655 10044 11667 10047
rect 12360 10044 12388 10084
rect 12710 10072 12716 10084
rect 12768 10072 12774 10124
rect 12897 10115 12955 10121
rect 12897 10081 12909 10115
rect 12943 10112 12955 10115
rect 15470 10112 15476 10124
rect 12943 10084 15476 10112
rect 12943 10081 12955 10084
rect 12897 10075 12955 10081
rect 15470 10072 15476 10084
rect 15528 10072 15534 10124
rect 22281 10115 22339 10121
rect 22281 10081 22293 10115
rect 22327 10112 22339 10115
rect 24578 10112 24584 10124
rect 22327 10084 24584 10112
rect 22327 10081 22339 10084
rect 22281 10075 22339 10081
rect 24578 10072 24584 10084
rect 24636 10072 24642 10124
rect 28353 10115 28411 10121
rect 28353 10081 28365 10115
rect 28399 10112 28411 10115
rect 29822 10112 29828 10124
rect 28399 10084 29828 10112
rect 28399 10081 28411 10084
rect 28353 10075 28411 10081
rect 29822 10072 29828 10084
rect 29880 10072 29886 10124
rect 29914 10072 29920 10124
rect 29972 10112 29978 10124
rect 30190 10112 30196 10124
rect 29972 10084 30196 10112
rect 29972 10072 29978 10084
rect 30190 10072 30196 10084
rect 30248 10112 30254 10124
rect 30285 10115 30343 10121
rect 30285 10112 30297 10115
rect 30248 10084 30297 10112
rect 30248 10072 30254 10084
rect 30285 10081 30297 10084
rect 30331 10081 30343 10115
rect 30285 10075 30343 10081
rect 30834 10072 30840 10124
rect 30892 10112 30898 10124
rect 32677 10115 32735 10121
rect 32677 10112 32689 10115
rect 30892 10084 32689 10112
rect 30892 10072 30898 10084
rect 32677 10081 32689 10084
rect 32723 10081 32735 10115
rect 32677 10075 32735 10081
rect 12621 10047 12679 10053
rect 12621 10044 12633 10047
rect 11655 10016 12296 10044
rect 12360 10016 12633 10044
rect 11655 10013 11667 10016
rect 11609 10007 11667 10013
rect 6362 9976 6368 9988
rect 6323 9948 6368 9976
rect 6362 9936 6368 9948
rect 6420 9936 6426 9988
rect 7650 9976 7656 9988
rect 7590 9948 7656 9976
rect 7650 9936 7656 9948
rect 7708 9936 7714 9988
rect 9401 9979 9459 9985
rect 9401 9976 9413 9979
rect 8588 9948 9413 9976
rect 7834 9908 7840 9920
rect 7795 9880 7840 9908
rect 7834 9868 7840 9880
rect 7892 9868 7898 9920
rect 8588 9917 8616 9948
rect 9401 9945 9413 9948
rect 9447 9945 9459 9979
rect 10778 9976 10784 9988
rect 10626 9948 10784 9976
rect 9401 9939 9459 9945
rect 10778 9936 10784 9948
rect 10836 9936 10842 9988
rect 8573 9911 8631 9917
rect 8573 9877 8585 9911
rect 8619 9877 8631 9911
rect 10870 9908 10876 9920
rect 10831 9880 10876 9908
rect 8573 9871 8631 9877
rect 10870 9868 10876 9880
rect 10928 9868 10934 9920
rect 12268 9917 12296 10016
rect 12621 10013 12633 10016
rect 12667 10044 12679 10047
rect 13906 10044 13912 10056
rect 12667 10016 13912 10044
rect 12667 10013 12679 10016
rect 12621 10007 12679 10013
rect 13906 10004 13912 10016
rect 13964 10004 13970 10056
rect 23658 10004 23664 10056
rect 23716 10004 23722 10056
rect 26418 10004 26424 10056
rect 26476 10044 26482 10056
rect 27525 10047 27583 10053
rect 27525 10044 27537 10047
rect 26476 10016 27537 10044
rect 26476 10004 26482 10016
rect 27525 10013 27537 10016
rect 27571 10013 27583 10047
rect 27525 10007 27583 10013
rect 28166 10004 28172 10056
rect 28224 10044 28230 10056
rect 29089 10047 29147 10053
rect 29089 10044 29101 10047
rect 28224 10016 29101 10044
rect 28224 10004 28230 10016
rect 29089 10013 29101 10016
rect 29135 10013 29147 10047
rect 29089 10007 29147 10013
rect 29454 10004 29460 10056
rect 29512 10044 29518 10056
rect 30101 10047 30159 10053
rect 30101 10044 30113 10047
rect 29512 10016 30113 10044
rect 29512 10004 29518 10016
rect 30101 10013 30113 10016
rect 30147 10013 30159 10047
rect 30101 10007 30159 10013
rect 31754 10004 31760 10056
rect 31812 10044 31818 10056
rect 33505 10047 33563 10053
rect 33505 10044 33517 10047
rect 31812 10016 33517 10044
rect 31812 10004 31818 10016
rect 33505 10013 33517 10016
rect 33551 10013 33563 10047
rect 33505 10007 33563 10013
rect 33594 10004 33600 10056
rect 33652 10044 33658 10056
rect 34149 10047 34207 10053
rect 34149 10044 34161 10047
rect 33652 10016 34161 10044
rect 33652 10004 33658 10016
rect 34149 10013 34161 10016
rect 34195 10013 34207 10047
rect 34149 10007 34207 10013
rect 22554 9976 22560 9988
rect 22515 9948 22560 9976
rect 22554 9936 22560 9948
rect 22612 9936 22618 9988
rect 24854 9976 24860 9988
rect 24815 9948 24860 9976
rect 24854 9936 24860 9948
rect 24912 9936 24918 9988
rect 25498 9936 25504 9988
rect 25556 9936 25562 9988
rect 27430 9936 27436 9988
rect 27488 9976 27494 9988
rect 31021 9979 31079 9985
rect 31021 9976 31033 9979
rect 27488 9948 31033 9976
rect 27488 9936 27494 9948
rect 31021 9945 31033 9948
rect 31067 9945 31079 9979
rect 31021 9939 31079 9945
rect 32493 9979 32551 9985
rect 32493 9945 32505 9979
rect 32539 9976 32551 9979
rect 33134 9976 33140 9988
rect 32539 9948 33140 9976
rect 32539 9945 32551 9948
rect 32493 9939 32551 9945
rect 33134 9936 33140 9948
rect 33192 9936 33198 9988
rect 12253 9911 12311 9917
rect 12253 9877 12265 9911
rect 12299 9877 12311 9911
rect 12253 9871 12311 9877
rect 30190 9868 30196 9920
rect 30248 9908 30254 9920
rect 32122 9908 32128 9920
rect 30248 9880 30293 9908
rect 32083 9880 32128 9908
rect 30248 9868 30254 9880
rect 32122 9868 32128 9880
rect 32180 9868 32186 9920
rect 32585 9911 32643 9917
rect 32585 9877 32597 9911
rect 32631 9908 32643 9911
rect 32950 9908 32956 9920
rect 32631 9880 32956 9908
rect 32631 9877 32643 9880
rect 32585 9871 32643 9877
rect 32950 9868 32956 9880
rect 33008 9868 33014 9920
rect 33410 9868 33416 9920
rect 33468 9908 33474 9920
rect 33965 9911 34023 9917
rect 33965 9908 33977 9911
rect 33468 9880 33977 9908
rect 33468 9868 33474 9880
rect 33965 9877 33977 9880
rect 34011 9877 34023 9911
rect 33965 9871 34023 9877
rect 1104 9818 37628 9840
rect 1104 9766 4874 9818
rect 4926 9766 4938 9818
rect 4990 9766 5002 9818
rect 5054 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 35594 9818
rect 35646 9766 35658 9818
rect 35710 9766 35722 9818
rect 35774 9766 35786 9818
rect 35838 9766 35850 9818
rect 35902 9766 37628 9818
rect 1104 9744 37628 9766
rect 8386 9664 8392 9716
rect 8444 9704 8450 9716
rect 8481 9707 8539 9713
rect 8481 9704 8493 9707
rect 8444 9676 8493 9704
rect 8444 9664 8450 9676
rect 8481 9673 8493 9676
rect 8527 9673 8539 9707
rect 8481 9667 8539 9673
rect 10045 9707 10103 9713
rect 10045 9673 10057 9707
rect 10091 9704 10103 9707
rect 10226 9704 10232 9716
rect 10091 9676 10232 9704
rect 10091 9673 10103 9676
rect 10045 9667 10103 9673
rect 10226 9664 10232 9676
rect 10284 9664 10290 9716
rect 12710 9664 12716 9716
rect 12768 9704 12774 9716
rect 13449 9707 13507 9713
rect 13449 9704 13461 9707
rect 12768 9676 13461 9704
rect 12768 9664 12774 9676
rect 13449 9673 13461 9676
rect 13495 9673 13507 9707
rect 13449 9667 13507 9673
rect 13906 9664 13912 9716
rect 13964 9704 13970 9716
rect 14369 9707 14427 9713
rect 14369 9704 14381 9707
rect 13964 9676 14381 9704
rect 13964 9664 13970 9676
rect 14369 9673 14381 9676
rect 14415 9673 14427 9707
rect 14369 9667 14427 9673
rect 23584 9676 23888 9704
rect 8849 9639 8907 9645
rect 8849 9636 8861 9639
rect 1780 9608 8861 9636
rect 1780 9577 1808 9608
rect 8849 9605 8861 9608
rect 8895 9636 8907 9639
rect 10137 9639 10195 9645
rect 10137 9636 10149 9639
rect 8895 9608 10149 9636
rect 8895 9605 8907 9608
rect 8849 9599 8907 9605
rect 10137 9605 10149 9608
rect 10183 9636 10195 9639
rect 10870 9636 10876 9648
rect 10183 9608 10876 9636
rect 10183 9605 10195 9608
rect 10137 9599 10195 9605
rect 10870 9596 10876 9608
rect 10928 9596 10934 9648
rect 12066 9596 12072 9648
rect 12124 9636 12130 9648
rect 12124 9608 12466 9636
rect 12124 9596 12130 9608
rect 22830 9596 22836 9648
rect 22888 9636 22894 9648
rect 23584 9636 23612 9676
rect 22888 9608 23612 9636
rect 22888 9596 22894 9608
rect 23658 9596 23664 9648
rect 23716 9636 23722 9648
rect 23753 9639 23811 9645
rect 23753 9636 23765 9639
rect 23716 9608 23765 9636
rect 23716 9596 23722 9608
rect 23753 9605 23765 9608
rect 23799 9605 23811 9639
rect 23753 9599 23811 9605
rect 23860 9636 23888 9676
rect 27706 9664 27712 9716
rect 27764 9704 27770 9716
rect 28721 9707 28779 9713
rect 28721 9704 28733 9707
rect 27764 9676 28733 9704
rect 27764 9664 27770 9676
rect 28721 9673 28733 9676
rect 28767 9673 28779 9707
rect 28721 9667 28779 9673
rect 28810 9664 28816 9716
rect 28868 9704 28874 9716
rect 28868 9676 28913 9704
rect 28868 9664 28874 9676
rect 25498 9636 25504 9648
rect 23860 9608 25084 9636
rect 25459 9608 25504 9636
rect 1765 9571 1823 9577
rect 1765 9537 1777 9571
rect 1811 9537 1823 9571
rect 1765 9531 1823 9537
rect 7098 9528 7104 9580
rect 7156 9568 7162 9580
rect 7377 9571 7435 9577
rect 7377 9568 7389 9571
rect 7156 9540 7389 9568
rect 7156 9528 7162 9540
rect 7377 9537 7389 9540
rect 7423 9537 7435 9571
rect 7377 9531 7435 9537
rect 7469 9571 7527 9577
rect 7469 9537 7481 9571
rect 7515 9568 7527 9571
rect 7834 9568 7840 9580
rect 7515 9540 7840 9568
rect 7515 9537 7527 9540
rect 7469 9531 7527 9537
rect 7834 9528 7840 9540
rect 7892 9528 7898 9580
rect 8294 9528 8300 9580
rect 8352 9568 8358 9580
rect 10962 9568 10968 9580
rect 8352 9540 9076 9568
rect 10923 9540 10968 9568
rect 8352 9528 8358 9540
rect 7650 9500 7656 9512
rect 7611 9472 7656 9500
rect 7650 9460 7656 9472
rect 7708 9460 7714 9512
rect 8202 9460 8208 9512
rect 8260 9500 8266 9512
rect 9048 9509 9076 9540
rect 10962 9528 10968 9540
rect 11020 9528 11026 9580
rect 11698 9568 11704 9580
rect 11659 9540 11704 9568
rect 11698 9528 11704 9540
rect 11756 9528 11762 9580
rect 14274 9568 14280 9580
rect 14235 9540 14280 9568
rect 14274 9528 14280 9540
rect 14332 9528 14338 9580
rect 23860 9577 23888 9608
rect 22649 9571 22707 9577
rect 22649 9537 22661 9571
rect 22695 9568 22707 9571
rect 23845 9571 23903 9577
rect 22695 9540 23796 9568
rect 22695 9537 22707 9540
rect 22649 9531 22707 9537
rect 8941 9503 8999 9509
rect 8941 9500 8953 9503
rect 8260 9472 8953 9500
rect 8260 9460 8266 9472
rect 8941 9469 8953 9472
rect 8987 9469 8999 9503
rect 8941 9463 8999 9469
rect 9033 9503 9091 9509
rect 9033 9469 9045 9503
rect 9079 9469 9091 9503
rect 9033 9463 9091 9469
rect 10229 9503 10287 9509
rect 10229 9469 10241 9503
rect 10275 9469 10287 9503
rect 11977 9503 12035 9509
rect 11977 9500 11989 9503
rect 10229 9463 10287 9469
rect 11164 9472 11989 9500
rect 6914 9392 6920 9444
rect 6972 9432 6978 9444
rect 7009 9435 7067 9441
rect 7009 9432 7021 9435
rect 6972 9404 7021 9432
rect 6972 9392 6978 9404
rect 7009 9401 7021 9404
rect 7055 9401 7067 9435
rect 7668 9432 7696 9460
rect 9766 9432 9772 9444
rect 7668 9404 9772 9432
rect 7009 9395 7067 9401
rect 9766 9392 9772 9404
rect 9824 9432 9830 9444
rect 10244 9432 10272 9463
rect 11164 9441 11192 9472
rect 11977 9469 11989 9472
rect 12023 9469 12035 9503
rect 11977 9463 12035 9469
rect 14553 9503 14611 9509
rect 14553 9469 14565 9503
rect 14599 9500 14611 9503
rect 15102 9500 15108 9512
rect 14599 9472 15108 9500
rect 14599 9469 14611 9472
rect 14553 9463 14611 9469
rect 15102 9460 15108 9472
rect 15160 9460 15166 9512
rect 22830 9500 22836 9512
rect 22791 9472 22836 9500
rect 22830 9460 22836 9472
rect 22888 9460 22894 9512
rect 23768 9500 23796 9540
rect 23845 9537 23857 9571
rect 23891 9537 23903 9571
rect 24946 9568 24952 9580
rect 24907 9540 24952 9568
rect 23845 9531 23903 9537
rect 24946 9528 24952 9540
rect 25004 9528 25010 9580
rect 25056 9568 25084 9608
rect 25498 9596 25504 9608
rect 25556 9596 25562 9648
rect 27614 9636 27620 9648
rect 27527 9608 27620 9636
rect 27614 9596 27620 9608
rect 27672 9636 27678 9648
rect 30190 9636 30196 9648
rect 27672 9608 30196 9636
rect 27672 9596 27678 9608
rect 30190 9596 30196 9608
rect 30248 9596 30254 9648
rect 30285 9639 30343 9645
rect 30285 9605 30297 9639
rect 30331 9636 30343 9639
rect 30374 9636 30380 9648
rect 30331 9608 30380 9636
rect 30331 9605 30343 9608
rect 30285 9599 30343 9605
rect 30374 9596 30380 9608
rect 30432 9596 30438 9648
rect 31662 9636 31668 9648
rect 31510 9608 31668 9636
rect 31662 9596 31668 9608
rect 31720 9596 31726 9648
rect 33137 9639 33195 9645
rect 33137 9605 33149 9639
rect 33183 9636 33195 9639
rect 33410 9636 33416 9648
rect 33183 9608 33416 9636
rect 33183 9605 33195 9608
rect 33137 9599 33195 9605
rect 33410 9596 33416 9608
rect 33468 9596 33474 9648
rect 33870 9596 33876 9648
rect 33928 9596 33934 9648
rect 25409 9571 25467 9577
rect 25409 9568 25421 9571
rect 25056 9540 25421 9568
rect 25409 9537 25421 9540
rect 25455 9568 25467 9571
rect 26053 9571 26111 9577
rect 26053 9568 26065 9571
rect 25455 9540 26065 9568
rect 25455 9537 25467 9540
rect 25409 9531 25467 9537
rect 26053 9537 26065 9540
rect 26099 9537 26111 9571
rect 26053 9531 26111 9537
rect 26234 9528 26240 9580
rect 26292 9528 26298 9580
rect 27525 9571 27583 9577
rect 27525 9537 27537 9571
rect 27571 9568 27583 9571
rect 27571 9540 28396 9568
rect 27571 9537 27583 9540
rect 27525 9531 27583 9537
rect 26252 9500 26280 9528
rect 27430 9500 27436 9512
rect 23768 9472 27436 9500
rect 27430 9460 27436 9472
rect 27488 9500 27494 9512
rect 27709 9503 27767 9509
rect 27709 9500 27721 9503
rect 27488 9472 27721 9500
rect 27488 9460 27494 9472
rect 27709 9469 27721 9472
rect 27755 9469 27767 9503
rect 27709 9463 27767 9469
rect 9824 9404 10272 9432
rect 11149 9435 11207 9441
rect 9824 9392 9830 9404
rect 11149 9401 11161 9435
rect 11195 9401 11207 9435
rect 11149 9395 11207 9401
rect 24765 9435 24823 9441
rect 24765 9401 24777 9435
rect 24811 9432 24823 9435
rect 24854 9432 24860 9444
rect 24811 9404 24860 9432
rect 24811 9401 24823 9404
rect 24765 9395 24823 9401
rect 24854 9392 24860 9404
rect 24912 9392 24918 9444
rect 28368 9441 28396 9540
rect 29822 9528 29828 9580
rect 29880 9568 29886 9580
rect 30009 9571 30067 9577
rect 30009 9568 30021 9571
rect 29880 9540 30021 9568
rect 29880 9528 29886 9540
rect 30009 9537 30021 9540
rect 30055 9537 30067 9571
rect 30009 9531 30067 9537
rect 28902 9460 28908 9512
rect 28960 9500 28966 9512
rect 28960 9472 29005 9500
rect 28960 9460 28966 9472
rect 28353 9435 28411 9441
rect 28353 9401 28365 9435
rect 28399 9401 28411 9435
rect 28353 9395 28411 9401
rect 1578 9364 1584 9376
rect 1539 9336 1584 9364
rect 1578 9324 1584 9336
rect 1636 9324 1642 9376
rect 9677 9367 9735 9373
rect 9677 9333 9689 9367
rect 9723 9364 9735 9367
rect 9858 9364 9864 9376
rect 9723 9336 9864 9364
rect 9723 9333 9735 9336
rect 9677 9327 9735 9333
rect 9858 9324 9864 9336
rect 9916 9324 9922 9376
rect 13906 9364 13912 9376
rect 13867 9336 13912 9364
rect 13906 9324 13912 9336
rect 13964 9324 13970 9376
rect 26050 9324 26056 9376
rect 26108 9364 26114 9376
rect 26145 9367 26203 9373
rect 26145 9364 26157 9367
rect 26108 9336 26157 9364
rect 26108 9324 26114 9336
rect 26145 9333 26157 9336
rect 26191 9333 26203 9367
rect 26145 9327 26203 9333
rect 26326 9324 26332 9376
rect 26384 9364 26390 9376
rect 27157 9367 27215 9373
rect 27157 9364 27169 9367
rect 26384 9336 27169 9364
rect 26384 9324 26390 9336
rect 27157 9333 27169 9336
rect 27203 9333 27215 9367
rect 30024 9364 30052 9531
rect 34422 9528 34428 9580
rect 34480 9568 34486 9580
rect 36725 9571 36783 9577
rect 36725 9568 36737 9571
rect 34480 9540 36737 9568
rect 34480 9528 34486 9540
rect 36725 9537 36737 9540
rect 36771 9537 36783 9571
rect 36725 9531 36783 9537
rect 31754 9500 31760 9512
rect 31312 9472 31760 9500
rect 31312 9364 31340 9472
rect 31754 9460 31760 9472
rect 31812 9500 31818 9512
rect 32861 9503 32919 9509
rect 32861 9500 32873 9503
rect 31812 9472 32873 9500
rect 31812 9460 31818 9472
rect 32861 9469 32873 9472
rect 32907 9469 32919 9503
rect 36906 9500 36912 9512
rect 32861 9463 32919 9469
rect 35866 9472 36912 9500
rect 30024 9336 31340 9364
rect 31757 9367 31815 9373
rect 27157 9327 27215 9333
rect 31757 9333 31769 9367
rect 31803 9364 31815 9367
rect 31846 9364 31852 9376
rect 31803 9336 31852 9364
rect 31803 9333 31815 9336
rect 31757 9327 31815 9333
rect 31846 9324 31852 9336
rect 31904 9324 31910 9376
rect 32950 9324 32956 9376
rect 33008 9364 33014 9376
rect 34609 9367 34667 9373
rect 34609 9364 34621 9367
rect 33008 9336 34621 9364
rect 33008 9324 33014 9336
rect 34609 9333 34621 9336
rect 34655 9364 34667 9367
rect 35866 9364 35894 9472
rect 36906 9460 36912 9472
rect 36964 9460 36970 9512
rect 36906 9364 36912 9376
rect 34655 9336 35894 9364
rect 36867 9336 36912 9364
rect 34655 9333 34667 9336
rect 34609 9327 34667 9333
rect 36906 9324 36912 9336
rect 36964 9324 36970 9376
rect 1104 9274 37628 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 37628 9274
rect 1104 9200 37628 9222
rect 7926 9120 7932 9172
rect 7984 9160 7990 9172
rect 10778 9160 10784 9172
rect 7984 9132 9996 9160
rect 10739 9132 10784 9160
rect 7984 9120 7990 9132
rect 8110 9052 8116 9104
rect 8168 9092 8174 9104
rect 8168 9064 9720 9092
rect 8168 9052 8174 9064
rect 6825 9027 6883 9033
rect 6825 8993 6837 9027
rect 6871 9024 6883 9027
rect 7190 9024 7196 9036
rect 6871 8996 7196 9024
rect 6871 8993 6883 8996
rect 6825 8987 6883 8993
rect 7190 8984 7196 8996
rect 7248 8984 7254 9036
rect 7650 8984 7656 9036
rect 7708 9024 7714 9036
rect 9692 9033 9720 9064
rect 8389 9027 8447 9033
rect 8389 9024 8401 9027
rect 7708 8996 8401 9024
rect 7708 8984 7714 8996
rect 8389 8993 8401 8996
rect 8435 8993 8447 9027
rect 8389 8987 8447 8993
rect 9677 9027 9735 9033
rect 9677 8993 9689 9027
rect 9723 8993 9735 9027
rect 9677 8987 9735 8993
rect 6181 8959 6239 8965
rect 6181 8925 6193 8959
rect 6227 8956 6239 8959
rect 7926 8956 7932 8968
rect 6227 8928 7932 8956
rect 6227 8925 6239 8928
rect 6181 8919 6239 8925
rect 7926 8916 7932 8928
rect 7984 8916 7990 8968
rect 8202 8956 8208 8968
rect 8163 8928 8208 8956
rect 8202 8916 8208 8928
rect 8260 8916 8266 8968
rect 9858 8956 9864 8968
rect 9819 8928 9864 8956
rect 9858 8916 9864 8928
rect 9916 8916 9922 8968
rect 9968 8956 9996 9132
rect 10778 9120 10784 9132
rect 10836 9120 10842 9172
rect 10962 9120 10968 9172
rect 11020 9160 11026 9172
rect 12069 9163 12127 9169
rect 12069 9160 12081 9163
rect 11020 9132 12081 9160
rect 11020 9120 11026 9132
rect 12069 9129 12081 9132
rect 12115 9129 12127 9163
rect 12069 9123 12127 9129
rect 26421 9163 26479 9169
rect 26421 9129 26433 9163
rect 26467 9160 26479 9163
rect 27614 9160 27620 9172
rect 26467 9132 27620 9160
rect 26467 9129 26479 9132
rect 26421 9123 26479 9129
rect 27614 9120 27620 9132
rect 27672 9120 27678 9172
rect 31386 9160 31392 9172
rect 31347 9132 31392 9160
rect 31386 9120 31392 9132
rect 31444 9120 31450 9172
rect 33321 9163 33379 9169
rect 33321 9129 33333 9163
rect 33367 9160 33379 9163
rect 33594 9160 33600 9172
rect 33367 9132 33600 9160
rect 33367 9129 33379 9132
rect 33321 9123 33379 9129
rect 33594 9120 33600 9132
rect 33652 9120 33658 9172
rect 33870 9120 33876 9172
rect 33928 9160 33934 9172
rect 33965 9163 34023 9169
rect 33965 9160 33977 9163
rect 33928 9132 33977 9160
rect 33928 9120 33934 9132
rect 33965 9129 33977 9132
rect 34011 9129 34023 9163
rect 33965 9123 34023 9129
rect 10229 9095 10287 9101
rect 10229 9061 10241 9095
rect 10275 9061 10287 9095
rect 14182 9092 14188 9104
rect 10229 9055 10287 9061
rect 12728 9064 14188 9092
rect 10244 9024 10272 9055
rect 12728 9033 12756 9064
rect 14182 9052 14188 9064
rect 14240 9052 14246 9104
rect 26234 9052 26240 9104
rect 26292 9092 26298 9104
rect 26292 9064 27016 9092
rect 26292 9052 26298 9064
rect 12713 9027 12771 9033
rect 10244 8996 11560 9024
rect 11532 8965 11560 8996
rect 12713 8993 12725 9027
rect 12759 8993 12771 9027
rect 13906 9024 13912 9036
rect 12713 8987 12771 8993
rect 13188 8996 13912 9024
rect 10873 8959 10931 8965
rect 10873 8956 10885 8959
rect 9968 8928 10885 8956
rect 10873 8925 10885 8928
rect 10919 8925 10931 8959
rect 10873 8919 10931 8925
rect 11517 8959 11575 8965
rect 11517 8925 11529 8959
rect 11563 8925 11575 8959
rect 11517 8919 11575 8925
rect 12437 8959 12495 8965
rect 12437 8925 12449 8959
rect 12483 8956 12495 8959
rect 13188 8956 13216 8996
rect 13906 8984 13912 8996
rect 13964 8984 13970 9036
rect 24578 8984 24584 9036
rect 24636 9024 24642 9036
rect 24673 9027 24731 9033
rect 24673 9024 24685 9027
rect 24636 8996 24685 9024
rect 24636 8984 24642 8996
rect 24673 8993 24685 8996
rect 24719 9024 24731 9027
rect 25682 9024 25688 9036
rect 24719 8996 25688 9024
rect 24719 8993 24731 8996
rect 24673 8987 24731 8993
rect 25682 8984 25688 8996
rect 25740 9024 25746 9036
rect 26881 9027 26939 9033
rect 26881 9024 26893 9027
rect 25740 8996 26893 9024
rect 25740 8984 25746 8996
rect 26881 8993 26893 8996
rect 26927 8993 26939 9027
rect 26988 9024 27016 9064
rect 28350 9024 28356 9036
rect 26988 8996 28356 9024
rect 26881 8987 26939 8993
rect 28350 8984 28356 8996
rect 28408 8984 28414 9036
rect 29178 8984 29184 9036
rect 29236 9024 29242 9036
rect 30561 9027 30619 9033
rect 30561 9024 30573 9027
rect 29236 8996 30573 9024
rect 29236 8984 29242 8996
rect 30561 8993 30573 8996
rect 30607 9024 30619 9027
rect 31110 9024 31116 9036
rect 30607 8996 31116 9024
rect 30607 8993 30619 8996
rect 30561 8987 30619 8993
rect 31110 8984 31116 8996
rect 31168 8984 31174 9036
rect 32030 9024 32036 9036
rect 31943 8996 32036 9024
rect 32030 8984 32036 8996
rect 32088 9024 32094 9036
rect 32490 9024 32496 9036
rect 32088 8996 32496 9024
rect 32088 8984 32094 8996
rect 32490 8984 32496 8996
rect 32548 8984 32554 9036
rect 32674 9024 32680 9036
rect 32635 8996 32680 9024
rect 32674 8984 32680 8996
rect 32732 9024 32738 9036
rect 33134 9024 33140 9036
rect 32732 8996 33140 9024
rect 32732 8984 32738 8996
rect 33134 8984 33140 8996
rect 33192 8984 33198 9036
rect 13538 8956 13544 8968
rect 12483 8928 13216 8956
rect 13499 8928 13544 8956
rect 12483 8925 12495 8928
rect 12437 8919 12495 8925
rect 13538 8916 13544 8928
rect 13596 8916 13602 8968
rect 13630 8916 13636 8968
rect 13688 8956 13694 8968
rect 14277 8959 14335 8965
rect 14277 8956 14289 8959
rect 13688 8928 14289 8956
rect 13688 8916 13694 8928
rect 14277 8925 14289 8928
rect 14323 8925 14335 8959
rect 14277 8919 14335 8925
rect 26050 8916 26056 8968
rect 26108 8916 26114 8968
rect 28368 8956 28396 8984
rect 29733 8959 29791 8965
rect 29733 8956 29745 8959
rect 28368 8928 29745 8956
rect 29733 8925 29745 8928
rect 29779 8925 29791 8959
rect 29733 8919 29791 8925
rect 31757 8959 31815 8965
rect 31757 8925 31769 8959
rect 31803 8956 31815 8959
rect 32122 8956 32128 8968
rect 31803 8928 32128 8956
rect 31803 8925 31815 8928
rect 31757 8919 31815 8925
rect 32122 8916 32128 8928
rect 32180 8916 32186 8968
rect 32950 8956 32956 8968
rect 32911 8928 32956 8956
rect 32950 8916 32956 8928
rect 33008 8916 33014 8968
rect 33778 8916 33784 8968
rect 33836 8956 33842 8968
rect 33873 8959 33931 8965
rect 33873 8956 33885 8959
rect 33836 8928 33885 8956
rect 33836 8916 33842 8928
rect 33873 8925 33885 8928
rect 33919 8956 33931 8959
rect 34790 8956 34796 8968
rect 33919 8928 34796 8956
rect 33919 8925 33931 8928
rect 33873 8919 33931 8925
rect 34790 8916 34796 8928
rect 34848 8916 34854 8968
rect 7009 8891 7067 8897
rect 7009 8857 7021 8891
rect 7055 8888 7067 8891
rect 8220 8888 8248 8916
rect 9769 8891 9827 8897
rect 9769 8888 9781 8891
rect 7055 8860 7880 8888
rect 8220 8860 9781 8888
rect 7055 8857 7067 8860
rect 7009 8851 7067 8857
rect 6086 8820 6092 8832
rect 6047 8792 6092 8820
rect 6086 8780 6092 8792
rect 6144 8780 6150 8832
rect 6917 8823 6975 8829
rect 6917 8789 6929 8823
rect 6963 8820 6975 8823
rect 7098 8820 7104 8832
rect 6963 8792 7104 8820
rect 6963 8789 6975 8792
rect 6917 8783 6975 8789
rect 7098 8780 7104 8792
rect 7156 8780 7162 8832
rect 7374 8820 7380 8832
rect 7335 8792 7380 8820
rect 7374 8780 7380 8792
rect 7432 8780 7438 8832
rect 7852 8829 7880 8860
rect 9769 8857 9781 8860
rect 9815 8857 9827 8891
rect 9769 8851 9827 8857
rect 12529 8891 12587 8897
rect 12529 8857 12541 8891
rect 12575 8888 12587 8891
rect 12710 8888 12716 8900
rect 12575 8860 12716 8888
rect 12575 8857 12587 8860
rect 12529 8851 12587 8857
rect 12710 8848 12716 8860
rect 12768 8848 12774 8900
rect 14550 8888 14556 8900
rect 14511 8860 14556 8888
rect 14550 8848 14556 8860
rect 14608 8848 14614 8900
rect 24946 8888 24952 8900
rect 14660 8860 15042 8888
rect 15856 8860 16574 8888
rect 24907 8860 24952 8888
rect 7837 8823 7895 8829
rect 7837 8789 7849 8823
rect 7883 8789 7895 8823
rect 7837 8783 7895 8789
rect 8018 8780 8024 8832
rect 8076 8820 8082 8832
rect 8297 8823 8355 8829
rect 8297 8820 8309 8823
rect 8076 8792 8309 8820
rect 8076 8780 8082 8792
rect 8297 8789 8309 8792
rect 8343 8789 8355 8823
rect 8297 8783 8355 8789
rect 10870 8780 10876 8832
rect 10928 8820 10934 8832
rect 11333 8823 11391 8829
rect 11333 8820 11345 8823
rect 10928 8792 11345 8820
rect 10928 8780 10934 8792
rect 11333 8789 11345 8792
rect 11379 8789 11391 8823
rect 11333 8783 11391 8789
rect 13633 8823 13691 8829
rect 13633 8789 13645 8823
rect 13679 8820 13691 8823
rect 14660 8820 14688 8860
rect 13679 8792 14688 8820
rect 13679 8789 13691 8792
rect 13633 8783 13691 8789
rect 15470 8780 15476 8832
rect 15528 8820 15534 8832
rect 15856 8820 15884 8860
rect 16022 8820 16028 8832
rect 15528 8792 15884 8820
rect 15983 8792 16028 8820
rect 15528 8780 15534 8792
rect 16022 8780 16028 8792
rect 16080 8780 16086 8832
rect 16546 8820 16574 8860
rect 24946 8848 24952 8860
rect 25004 8848 25010 8900
rect 27154 8888 27160 8900
rect 27115 8860 27160 8888
rect 27154 8848 27160 8860
rect 27212 8848 27218 8900
rect 27614 8848 27620 8900
rect 27672 8848 27678 8900
rect 31846 8888 31852 8900
rect 31759 8860 31852 8888
rect 31846 8848 31852 8860
rect 31904 8888 31910 8900
rect 32861 8891 32919 8897
rect 32861 8888 32873 8891
rect 31904 8860 32873 8888
rect 31904 8848 31910 8860
rect 32861 8857 32873 8860
rect 32907 8888 32919 8891
rect 33594 8888 33600 8900
rect 32907 8860 33600 8888
rect 32907 8857 32919 8860
rect 32861 8851 32919 8857
rect 33594 8848 33600 8860
rect 33652 8848 33658 8900
rect 22278 8820 22284 8832
rect 16546 8792 22284 8820
rect 22278 8780 22284 8792
rect 22336 8820 22342 8832
rect 22830 8820 22836 8832
rect 22336 8792 22836 8820
rect 22336 8780 22342 8792
rect 22830 8780 22836 8792
rect 22888 8780 22894 8832
rect 28626 8820 28632 8832
rect 28587 8792 28632 8820
rect 28626 8780 28632 8792
rect 28684 8780 28690 8832
rect 1104 8730 37628 8752
rect 1104 8678 4874 8730
rect 4926 8678 4938 8730
rect 4990 8678 5002 8730
rect 5054 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 35594 8730
rect 35646 8678 35658 8730
rect 35710 8678 35722 8730
rect 35774 8678 35786 8730
rect 35838 8678 35850 8730
rect 35902 8678 37628 8730
rect 1104 8656 37628 8678
rect 8202 8576 8208 8628
rect 8260 8616 8266 8628
rect 9401 8619 9459 8625
rect 9401 8616 9413 8619
rect 8260 8588 9413 8616
rect 8260 8576 8266 8588
rect 9401 8585 9413 8588
rect 9447 8585 9459 8619
rect 12066 8616 12072 8628
rect 12027 8588 12072 8616
rect 9401 8579 9459 8585
rect 12066 8576 12072 8588
rect 12124 8576 12130 8628
rect 13633 8619 13691 8625
rect 13633 8585 13645 8619
rect 13679 8616 13691 8619
rect 14550 8616 14556 8628
rect 13679 8588 14556 8616
rect 13679 8585 13691 8588
rect 13633 8579 13691 8585
rect 14550 8576 14556 8588
rect 14608 8576 14614 8628
rect 15562 8576 15568 8628
rect 15620 8616 15626 8628
rect 15841 8619 15899 8625
rect 15841 8616 15853 8619
rect 15620 8588 15853 8616
rect 15620 8576 15626 8588
rect 15841 8585 15853 8588
rect 15887 8616 15899 8619
rect 26418 8616 26424 8628
rect 15887 8588 18644 8616
rect 15887 8585 15899 8588
rect 15841 8579 15899 8585
rect 6086 8508 6092 8560
rect 6144 8548 6150 8560
rect 6144 8520 6854 8548
rect 6144 8508 6150 8520
rect 10410 8508 10416 8560
rect 10468 8508 10474 8560
rect 10870 8548 10876 8560
rect 10831 8520 10876 8548
rect 10870 8508 10876 8520
rect 10928 8508 10934 8560
rect 12434 8548 12440 8560
rect 11992 8520 12440 8548
rect 5810 8480 5816 8492
rect 5771 8452 5816 8480
rect 5810 8440 5816 8452
rect 5868 8440 5874 8492
rect 11992 8489 12020 8520
rect 12434 8508 12440 8520
rect 12492 8548 12498 8560
rect 13538 8548 13544 8560
rect 12492 8520 13544 8548
rect 12492 8508 12498 8520
rect 13538 8508 13544 8520
rect 13596 8508 13602 8560
rect 14274 8508 14280 8560
rect 14332 8548 14338 8560
rect 15749 8551 15807 8557
rect 15749 8548 15761 8551
rect 14332 8520 15761 8548
rect 14332 8508 14338 8520
rect 11977 8483 12035 8489
rect 11977 8449 11989 8483
rect 12023 8449 12035 8483
rect 11977 8443 12035 8449
rect 13449 8483 13507 8489
rect 13449 8449 13461 8483
rect 13495 8480 13507 8483
rect 14458 8480 14464 8492
rect 13495 8452 14136 8480
rect 14419 8452 14464 8480
rect 13495 8449 13507 8452
rect 13449 8443 13507 8449
rect 8021 8415 8079 8421
rect 8021 8412 8033 8415
rect 6012 8384 8033 8412
rect 6012 8353 6040 8384
rect 8021 8381 8033 8384
rect 8067 8381 8079 8415
rect 8021 8375 8079 8381
rect 8297 8415 8355 8421
rect 8297 8381 8309 8415
rect 8343 8412 8355 8415
rect 9214 8412 9220 8424
rect 8343 8384 9220 8412
rect 8343 8381 8355 8384
rect 8297 8375 8355 8381
rect 9214 8372 9220 8384
rect 9272 8372 9278 8424
rect 11149 8415 11207 8421
rect 11149 8381 11161 8415
rect 11195 8412 11207 8415
rect 11790 8412 11796 8424
rect 11195 8384 11796 8412
rect 11195 8381 11207 8384
rect 11149 8375 11207 8381
rect 11790 8372 11796 8384
rect 11848 8412 11854 8424
rect 13630 8412 13636 8424
rect 11848 8384 13636 8412
rect 11848 8372 11854 8384
rect 13630 8372 13636 8384
rect 13688 8372 13694 8424
rect 5997 8347 6055 8353
rect 5997 8313 6009 8347
rect 6043 8313 6055 8347
rect 5997 8307 6055 8313
rect 6549 8347 6607 8353
rect 6549 8313 6561 8347
rect 6595 8344 6607 8347
rect 7006 8344 7012 8356
rect 6595 8316 7012 8344
rect 6595 8313 6607 8316
rect 6549 8307 6607 8313
rect 7006 8304 7012 8316
rect 7064 8304 7070 8356
rect 14108 8353 14136 8452
rect 14458 8440 14464 8452
rect 14516 8440 14522 8492
rect 14568 8489 14596 8520
rect 15749 8517 15761 8520
rect 15795 8548 15807 8551
rect 16022 8548 16028 8560
rect 15795 8520 16028 8548
rect 15795 8517 15807 8520
rect 15749 8511 15807 8517
rect 16022 8508 16028 8520
rect 16080 8508 16086 8560
rect 18138 8508 18144 8560
rect 18196 8508 18202 8560
rect 14553 8483 14611 8489
rect 14553 8449 14565 8483
rect 14599 8449 14611 8483
rect 14553 8443 14611 8449
rect 14645 8415 14703 8421
rect 14645 8381 14657 8415
rect 14691 8381 14703 8415
rect 14645 8375 14703 8381
rect 14093 8347 14151 8353
rect 14093 8313 14105 8347
rect 14139 8313 14151 8347
rect 14093 8307 14151 8313
rect 14182 8304 14188 8356
rect 14240 8344 14246 8356
rect 14550 8344 14556 8356
rect 14240 8316 14556 8344
rect 14240 8304 14246 8316
rect 14550 8304 14556 8316
rect 14608 8344 14614 8356
rect 14660 8344 14688 8375
rect 15470 8372 15476 8424
rect 15528 8412 15534 8424
rect 15565 8415 15623 8421
rect 15565 8412 15577 8415
rect 15528 8384 15577 8412
rect 15528 8372 15534 8384
rect 15565 8381 15577 8384
rect 15611 8381 15623 8415
rect 15565 8375 15623 8381
rect 16022 8372 16028 8424
rect 16080 8412 16086 8424
rect 16853 8415 16911 8421
rect 16853 8412 16865 8415
rect 16080 8384 16865 8412
rect 16080 8372 16086 8384
rect 16853 8381 16865 8384
rect 16899 8381 16911 8415
rect 17126 8412 17132 8424
rect 17087 8384 17132 8412
rect 16853 8375 16911 8381
rect 17126 8372 17132 8384
rect 17184 8372 17190 8424
rect 18616 8353 18644 8588
rect 26206 8588 26424 8616
rect 25041 8551 25099 8557
rect 25041 8517 25053 8551
rect 25087 8548 25099 8551
rect 26206 8548 26234 8588
rect 26418 8576 26424 8588
rect 26476 8576 26482 8628
rect 26513 8619 26571 8625
rect 26513 8585 26525 8619
rect 26559 8616 26571 8619
rect 27614 8616 27620 8628
rect 26559 8588 27620 8616
rect 26559 8585 26571 8588
rect 26513 8579 26571 8585
rect 27614 8576 27620 8588
rect 27672 8576 27678 8628
rect 27801 8619 27859 8625
rect 27801 8585 27813 8619
rect 27847 8616 27859 8619
rect 28626 8616 28632 8628
rect 27847 8588 28632 8616
rect 27847 8585 27859 8588
rect 27801 8579 27859 8585
rect 28626 8576 28632 8588
rect 28684 8576 28690 8628
rect 30469 8619 30527 8625
rect 30469 8585 30481 8619
rect 30515 8616 30527 8619
rect 30650 8616 30656 8628
rect 30515 8588 30656 8616
rect 30515 8585 30527 8588
rect 30469 8579 30527 8585
rect 30650 8576 30656 8588
rect 30708 8576 30714 8628
rect 31662 8616 31668 8628
rect 31623 8588 31668 8616
rect 31662 8576 31668 8588
rect 31720 8576 31726 8628
rect 32677 8619 32735 8625
rect 32677 8585 32689 8619
rect 32723 8616 32735 8619
rect 33505 8619 33563 8625
rect 33505 8616 33517 8619
rect 32723 8588 33517 8616
rect 32723 8585 32735 8588
rect 32677 8579 32735 8585
rect 33505 8585 33517 8588
rect 33551 8585 33563 8619
rect 33505 8579 33563 8585
rect 33594 8576 33600 8628
rect 33652 8616 33658 8628
rect 33873 8619 33931 8625
rect 33873 8616 33885 8619
rect 33652 8588 33885 8616
rect 33652 8576 33658 8588
rect 33873 8585 33885 8588
rect 33919 8585 33931 8619
rect 33873 8579 33931 8585
rect 33965 8619 34023 8625
rect 33965 8585 33977 8619
rect 34011 8616 34023 8619
rect 34330 8616 34336 8628
rect 34011 8588 34336 8616
rect 34011 8585 34023 8588
rect 33965 8579 34023 8585
rect 34330 8576 34336 8588
rect 34388 8576 34394 8628
rect 30282 8548 30288 8560
rect 25087 8520 26234 8548
rect 26344 8520 28764 8548
rect 30222 8520 30288 8548
rect 25087 8517 25099 8520
rect 25041 8511 25099 8517
rect 25682 8440 25688 8492
rect 25740 8480 25746 8492
rect 25777 8483 25835 8489
rect 25777 8480 25789 8483
rect 25740 8452 25789 8480
rect 25740 8440 25746 8452
rect 25777 8449 25789 8452
rect 25823 8480 25835 8483
rect 26050 8480 26056 8492
rect 25823 8452 26056 8480
rect 25823 8449 25835 8452
rect 25777 8443 25835 8449
rect 26050 8440 26056 8452
rect 26108 8480 26114 8492
rect 26344 8480 26372 8520
rect 26108 8452 26372 8480
rect 26421 8483 26479 8489
rect 26108 8440 26114 8452
rect 26421 8449 26433 8483
rect 26467 8480 26479 8483
rect 27798 8480 27804 8492
rect 26467 8452 27804 8480
rect 26467 8449 26479 8452
rect 26421 8443 26479 8449
rect 27798 8440 27804 8452
rect 27856 8440 27862 8492
rect 27893 8483 27951 8489
rect 27893 8449 27905 8483
rect 27939 8480 27951 8483
rect 27982 8480 27988 8492
rect 27939 8452 27988 8480
rect 27939 8449 27951 8452
rect 27893 8443 27951 8449
rect 27982 8440 27988 8452
rect 28040 8440 28046 8492
rect 28736 8489 28764 8520
rect 30282 8508 30288 8520
rect 30340 8508 30346 8560
rect 30834 8508 30840 8560
rect 30892 8548 30898 8560
rect 30892 8520 34100 8548
rect 30892 8508 30898 8520
rect 28721 8483 28779 8489
rect 28721 8449 28733 8483
rect 28767 8449 28779 8483
rect 31110 8480 31116 8492
rect 31071 8452 31116 8480
rect 28721 8443 28779 8449
rect 31110 8440 31116 8452
rect 31168 8440 31174 8492
rect 31757 8483 31815 8489
rect 31757 8449 31769 8483
rect 31803 8480 31815 8483
rect 32858 8480 32864 8492
rect 31803 8452 32864 8480
rect 31803 8449 31815 8452
rect 31757 8443 31815 8449
rect 32858 8440 32864 8452
rect 32916 8440 32922 8492
rect 27709 8415 27767 8421
rect 27709 8381 27721 8415
rect 27755 8381 27767 8415
rect 27709 8375 27767 8381
rect 28997 8415 29055 8421
rect 28997 8381 29009 8415
rect 29043 8412 29055 8415
rect 32490 8412 32496 8424
rect 29043 8384 30972 8412
rect 32451 8384 32496 8412
rect 29043 8381 29055 8384
rect 28997 8375 29055 8381
rect 14608 8316 14688 8344
rect 18601 8347 18659 8353
rect 14608 8304 14614 8316
rect 18601 8313 18613 8347
rect 18647 8344 18659 8347
rect 21450 8344 21456 8356
rect 18647 8316 21456 8344
rect 18647 8313 18659 8316
rect 18601 8307 18659 8313
rect 21450 8304 21456 8316
rect 21508 8304 21514 8356
rect 27724 8344 27752 8375
rect 28718 8344 28724 8356
rect 27724 8316 28724 8344
rect 28718 8304 28724 8316
rect 28776 8304 28782 8356
rect 30944 8353 30972 8384
rect 32490 8372 32496 8384
rect 32548 8372 32554 8424
rect 32585 8415 32643 8421
rect 32585 8381 32597 8415
rect 32631 8412 32643 8415
rect 32766 8412 32772 8424
rect 32631 8384 32772 8412
rect 32631 8381 32643 8384
rect 32585 8375 32643 8381
rect 32766 8372 32772 8384
rect 32824 8372 32830 8424
rect 34072 8421 34100 8520
rect 34790 8440 34796 8492
rect 34848 8480 34854 8492
rect 34885 8483 34943 8489
rect 34885 8480 34897 8483
rect 34848 8452 34897 8480
rect 34848 8440 34854 8452
rect 34885 8449 34897 8452
rect 34931 8449 34943 8483
rect 34885 8443 34943 8449
rect 34057 8415 34115 8421
rect 34057 8381 34069 8415
rect 34103 8381 34115 8415
rect 34057 8375 34115 8381
rect 30929 8347 30987 8353
rect 30929 8313 30941 8347
rect 30975 8313 30987 8347
rect 30929 8307 30987 8313
rect 33045 8347 33103 8353
rect 33045 8313 33057 8347
rect 33091 8344 33103 8347
rect 34606 8344 34612 8356
rect 33091 8316 34612 8344
rect 33091 8313 33103 8316
rect 33045 8307 33103 8313
rect 34606 8304 34612 8316
rect 34664 8304 34670 8356
rect 34790 8344 34796 8356
rect 34751 8316 34796 8344
rect 34790 8304 34796 8316
rect 34848 8304 34854 8356
rect 16209 8279 16267 8285
rect 16209 8245 16221 8279
rect 16255 8276 16267 8279
rect 16298 8276 16304 8288
rect 16255 8248 16304 8276
rect 16255 8245 16267 8248
rect 16209 8239 16267 8245
rect 16298 8236 16304 8248
rect 16356 8236 16362 8288
rect 28261 8279 28319 8285
rect 28261 8245 28273 8279
rect 28307 8276 28319 8279
rect 28810 8276 28816 8288
rect 28307 8248 28816 8276
rect 28307 8245 28319 8248
rect 28261 8239 28319 8245
rect 28810 8236 28816 8248
rect 28868 8236 28874 8288
rect 1104 8186 37628 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 37628 8186
rect 1104 8112 37628 8134
rect 5810 8032 5816 8084
rect 5868 8072 5874 8084
rect 6733 8075 6791 8081
rect 6733 8072 6745 8075
rect 5868 8044 6745 8072
rect 5868 8032 5874 8044
rect 6733 8041 6745 8044
rect 6779 8041 6791 8075
rect 6733 8035 6791 8041
rect 10410 8032 10416 8084
rect 10468 8072 10474 8084
rect 10689 8075 10747 8081
rect 10689 8072 10701 8075
rect 10468 8044 10701 8072
rect 10468 8032 10474 8044
rect 10689 8041 10701 8044
rect 10735 8041 10747 8075
rect 10689 8035 10747 8041
rect 14458 8032 14464 8084
rect 14516 8072 14522 8084
rect 15105 8075 15163 8081
rect 15105 8072 15117 8075
rect 14516 8044 15117 8072
rect 14516 8032 14522 8044
rect 15105 8041 15117 8044
rect 15151 8041 15163 8075
rect 15105 8035 15163 8041
rect 16485 8075 16543 8081
rect 16485 8041 16497 8075
rect 16531 8072 16543 8075
rect 17126 8072 17132 8084
rect 16531 8044 17132 8072
rect 16531 8041 16543 8044
rect 16485 8035 16543 8041
rect 17126 8032 17132 8044
rect 17184 8032 17190 8084
rect 17313 8075 17371 8081
rect 17313 8041 17325 8075
rect 17359 8072 17371 8075
rect 18138 8072 18144 8084
rect 17359 8044 18144 8072
rect 17359 8041 17371 8044
rect 17313 8035 17371 8041
rect 18138 8032 18144 8044
rect 18196 8032 18202 8084
rect 24946 8032 24952 8084
rect 25004 8072 25010 8084
rect 25317 8075 25375 8081
rect 25317 8072 25329 8075
rect 25004 8044 25329 8072
rect 25004 8032 25010 8044
rect 25317 8041 25329 8044
rect 25363 8041 25375 8075
rect 27154 8072 27160 8084
rect 27115 8044 27160 8072
rect 25317 8035 25375 8041
rect 27154 8032 27160 8044
rect 27212 8032 27218 8084
rect 30469 8075 30527 8081
rect 30469 8041 30481 8075
rect 30515 8072 30527 8075
rect 31110 8072 31116 8084
rect 30515 8044 31116 8072
rect 30515 8041 30527 8044
rect 30469 8035 30527 8041
rect 31110 8032 31116 8044
rect 31168 8032 31174 8084
rect 31284 8075 31342 8081
rect 31284 8041 31296 8075
rect 31330 8072 31342 8075
rect 34885 8075 34943 8081
rect 34885 8072 34897 8075
rect 31330 8044 34897 8072
rect 31330 8041 31342 8044
rect 31284 8035 31342 8041
rect 34885 8041 34897 8044
rect 34931 8041 34943 8075
rect 34885 8035 34943 8041
rect 15194 7964 15200 8016
rect 15252 8004 15258 8016
rect 15378 8004 15384 8016
rect 15252 7976 15384 8004
rect 15252 7964 15258 7976
rect 15378 7964 15384 7976
rect 15436 8004 15442 8016
rect 28353 8007 28411 8013
rect 15436 7976 15700 8004
rect 15436 7964 15442 7976
rect 7098 7896 7104 7948
rect 7156 7936 7162 7948
rect 7193 7939 7251 7945
rect 7193 7936 7205 7939
rect 7156 7908 7205 7936
rect 7156 7896 7162 7908
rect 7193 7905 7205 7908
rect 7239 7905 7251 7939
rect 7193 7899 7251 7905
rect 7285 7939 7343 7945
rect 7285 7905 7297 7939
rect 7331 7936 7343 7939
rect 8294 7936 8300 7948
rect 7331 7908 8300 7936
rect 7331 7905 7343 7908
rect 7285 7899 7343 7905
rect 8294 7896 8300 7908
rect 8352 7896 8358 7948
rect 13630 7936 13636 7948
rect 13591 7908 13636 7936
rect 13630 7896 13636 7908
rect 13688 7896 13694 7948
rect 15562 7936 15568 7948
rect 15523 7908 15568 7936
rect 15562 7896 15568 7908
rect 15620 7896 15626 7948
rect 15672 7945 15700 7976
rect 28353 7973 28365 8007
rect 28399 7973 28411 8007
rect 30558 8004 30564 8016
rect 28353 7967 28411 7973
rect 28920 7976 30564 8004
rect 15657 7939 15715 7945
rect 15657 7905 15669 7939
rect 15703 7905 15715 7939
rect 15657 7899 15715 7905
rect 7374 7828 7380 7880
rect 7432 7868 7438 7880
rect 7929 7871 7987 7877
rect 7929 7868 7941 7871
rect 7432 7840 7941 7868
rect 7432 7828 7438 7840
rect 7929 7837 7941 7840
rect 7975 7837 7987 7871
rect 7929 7831 7987 7837
rect 9309 7871 9367 7877
rect 9309 7837 9321 7871
rect 9355 7868 9367 7871
rect 10781 7871 10839 7877
rect 10781 7868 10793 7871
rect 9355 7840 10793 7868
rect 9355 7837 9367 7840
rect 9309 7831 9367 7837
rect 10781 7837 10793 7840
rect 10827 7868 10839 7871
rect 12434 7868 12440 7880
rect 10827 7840 12440 7868
rect 10827 7837 10839 7840
rect 10781 7831 10839 7837
rect 12434 7828 12440 7840
rect 12492 7828 12498 7880
rect 13538 7828 13544 7880
rect 13596 7868 13602 7880
rect 14277 7871 14335 7877
rect 14277 7868 14289 7871
rect 13596 7840 14289 7868
rect 13596 7828 13602 7840
rect 14277 7837 14289 7840
rect 14323 7837 14335 7871
rect 16298 7868 16304 7880
rect 16259 7840 16304 7868
rect 14277 7831 14335 7837
rect 16298 7828 16304 7840
rect 16356 7828 16362 7880
rect 17218 7868 17224 7880
rect 17179 7840 17224 7868
rect 17218 7828 17224 7840
rect 17276 7828 17282 7880
rect 25501 7871 25559 7877
rect 25501 7837 25513 7871
rect 25547 7868 25559 7871
rect 26326 7868 26332 7880
rect 25547 7840 26332 7868
rect 25547 7837 25559 7840
rect 25501 7831 25559 7837
rect 26326 7828 26332 7840
rect 26384 7828 26390 7880
rect 27341 7871 27399 7877
rect 27341 7837 27353 7871
rect 27387 7868 27399 7871
rect 28368 7868 28396 7967
rect 28920 7948 28948 7976
rect 30558 7964 30564 7976
rect 30616 8004 30622 8016
rect 30926 8004 30932 8016
rect 30616 7976 30932 8004
rect 30616 7964 30622 7976
rect 30926 7964 30932 7976
rect 30984 7964 30990 8016
rect 28902 7936 28908 7948
rect 28815 7908 28908 7936
rect 28902 7896 28908 7908
rect 28960 7896 28966 7948
rect 29914 7936 29920 7948
rect 29875 7908 29920 7936
rect 29914 7896 29920 7908
rect 29972 7896 29978 7948
rect 30009 7939 30067 7945
rect 30009 7905 30021 7939
rect 30055 7936 30067 7939
rect 30650 7936 30656 7948
rect 30055 7908 30656 7936
rect 30055 7905 30067 7908
rect 30009 7899 30067 7905
rect 27387 7840 28396 7868
rect 27387 7837 27399 7840
rect 27341 7831 27399 7837
rect 28626 7828 28632 7880
rect 28684 7868 28690 7880
rect 28721 7871 28779 7877
rect 28721 7868 28733 7871
rect 28684 7840 28733 7868
rect 28684 7828 28690 7840
rect 28721 7837 28733 7840
rect 28767 7837 28779 7871
rect 28721 7831 28779 7837
rect 28810 7828 28816 7880
rect 28868 7868 28874 7880
rect 30101 7871 30159 7877
rect 30101 7868 30113 7871
rect 28868 7840 30113 7868
rect 28868 7828 28874 7840
rect 30101 7837 30113 7840
rect 30147 7837 30159 7871
rect 30101 7831 30159 7837
rect 7006 7760 7012 7812
rect 7064 7800 7070 7812
rect 7101 7803 7159 7809
rect 7101 7800 7113 7803
rect 7064 7772 7113 7800
rect 7064 7760 7070 7772
rect 7101 7769 7113 7772
rect 7147 7800 7159 7803
rect 8018 7800 8024 7812
rect 7147 7772 8024 7800
rect 7147 7769 7159 7772
rect 7101 7763 7159 7769
rect 8018 7760 8024 7772
rect 8076 7760 8082 7812
rect 12618 7760 12624 7812
rect 12676 7800 12682 7812
rect 12805 7803 12863 7809
rect 12805 7800 12817 7803
rect 12676 7772 12817 7800
rect 12676 7760 12682 7772
rect 12805 7769 12817 7772
rect 12851 7800 12863 7803
rect 16206 7800 16212 7812
rect 12851 7772 16212 7800
rect 12851 7769 12863 7772
rect 12805 7763 12863 7769
rect 16206 7760 16212 7772
rect 16264 7760 16270 7812
rect 8113 7735 8171 7741
rect 8113 7701 8125 7735
rect 8159 7732 8171 7735
rect 8938 7732 8944 7744
rect 8159 7704 8944 7732
rect 8159 7701 8171 7704
rect 8113 7695 8171 7701
rect 8938 7692 8944 7704
rect 8996 7692 9002 7744
rect 9030 7692 9036 7744
rect 9088 7732 9094 7744
rect 9217 7735 9275 7741
rect 9217 7732 9229 7735
rect 9088 7704 9229 7732
rect 9088 7692 9094 7704
rect 9217 7701 9229 7704
rect 9263 7701 9275 7735
rect 14366 7732 14372 7744
rect 14327 7704 14372 7732
rect 9217 7695 9275 7701
rect 14366 7692 14372 7704
rect 14424 7692 14430 7744
rect 15470 7732 15476 7744
rect 15431 7704 15476 7732
rect 15470 7692 15476 7704
rect 15528 7692 15534 7744
rect 28813 7735 28871 7741
rect 28813 7701 28825 7735
rect 28859 7732 28871 7735
rect 30208 7732 30236 7908
rect 30650 7896 30656 7908
rect 30708 7896 30714 7948
rect 31021 7939 31079 7945
rect 31021 7905 31033 7939
rect 31067 7936 31079 7939
rect 31754 7936 31760 7948
rect 31067 7908 31760 7936
rect 31067 7905 31079 7908
rect 31021 7899 31079 7905
rect 31754 7896 31760 7908
rect 31812 7896 31818 7948
rect 33134 7896 33140 7948
rect 33192 7936 33198 7948
rect 33321 7939 33379 7945
rect 33321 7936 33333 7939
rect 33192 7908 33333 7936
rect 33192 7896 33198 7908
rect 33321 7905 33333 7908
rect 33367 7905 33379 7939
rect 33321 7899 33379 7905
rect 33597 7871 33655 7877
rect 33597 7837 33609 7871
rect 33643 7868 33655 7871
rect 34330 7868 34336 7880
rect 33643 7840 34336 7868
rect 33643 7837 33655 7840
rect 33597 7831 33655 7837
rect 34330 7828 34336 7840
rect 34388 7828 34394 7880
rect 34606 7828 34612 7880
rect 34664 7868 34670 7880
rect 35069 7871 35127 7877
rect 35069 7868 35081 7871
rect 34664 7840 35081 7868
rect 34664 7828 34670 7840
rect 35069 7837 35081 7840
rect 35115 7837 35127 7871
rect 35069 7831 35127 7837
rect 32950 7800 32956 7812
rect 32522 7772 32956 7800
rect 32950 7760 32956 7772
rect 33008 7760 33014 7812
rect 32766 7732 32772 7744
rect 28859 7704 30236 7732
rect 32727 7704 32772 7732
rect 28859 7701 28871 7704
rect 28813 7695 28871 7701
rect 32766 7692 32772 7704
rect 32824 7732 32830 7744
rect 33505 7735 33563 7741
rect 33505 7732 33517 7735
rect 32824 7704 33517 7732
rect 32824 7692 32830 7704
rect 33505 7701 33517 7704
rect 33551 7701 33563 7735
rect 33505 7695 33563 7701
rect 33965 7735 34023 7741
rect 33965 7701 33977 7735
rect 34011 7732 34023 7735
rect 34146 7732 34152 7744
rect 34011 7704 34152 7732
rect 34011 7701 34023 7704
rect 33965 7695 34023 7701
rect 34146 7692 34152 7704
rect 34204 7692 34210 7744
rect 1104 7642 37628 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 35594 7642
rect 35646 7590 35658 7642
rect 35710 7590 35722 7642
rect 35774 7590 35786 7642
rect 35838 7590 35850 7642
rect 35902 7590 37628 7642
rect 1104 7568 37628 7590
rect 7098 7488 7104 7540
rect 7156 7528 7162 7540
rect 7469 7531 7527 7537
rect 7469 7528 7481 7531
rect 7156 7500 7481 7528
rect 7156 7488 7162 7500
rect 7469 7497 7481 7500
rect 7515 7497 7527 7531
rect 9030 7528 9036 7540
rect 7469 7491 7527 7497
rect 8588 7500 9036 7528
rect 8588 7460 8616 7500
rect 9030 7488 9036 7500
rect 9088 7488 9094 7540
rect 15749 7531 15807 7537
rect 15749 7528 15761 7531
rect 15028 7500 15761 7528
rect 8938 7460 8944 7472
rect 8510 7432 8616 7460
rect 8899 7432 8944 7460
rect 8938 7420 8944 7432
rect 8996 7420 9002 7472
rect 14366 7420 14372 7472
rect 14424 7420 14430 7472
rect 15028 7469 15056 7500
rect 15749 7497 15761 7500
rect 15795 7497 15807 7531
rect 15749 7491 15807 7497
rect 28000 7500 30144 7528
rect 15013 7463 15071 7469
rect 15013 7429 15025 7463
rect 15059 7429 15071 7463
rect 15013 7423 15071 7429
rect 9214 7352 9220 7404
rect 9272 7392 9278 7404
rect 11790 7392 11796 7404
rect 9272 7364 11796 7392
rect 9272 7352 9278 7364
rect 11790 7352 11796 7364
rect 11848 7352 11854 7404
rect 12342 7392 12348 7404
rect 12303 7364 12348 7392
rect 12342 7352 12348 7364
rect 12400 7352 12406 7404
rect 12434 7352 12440 7404
rect 12492 7392 12498 7404
rect 12805 7395 12863 7401
rect 12805 7392 12817 7395
rect 12492 7364 12817 7392
rect 12492 7352 12498 7364
rect 12805 7361 12817 7364
rect 12851 7361 12863 7395
rect 15930 7392 15936 7404
rect 15891 7364 15936 7392
rect 12805 7355 12863 7361
rect 15930 7352 15936 7364
rect 15988 7352 15994 7404
rect 27338 7392 27344 7404
rect 27299 7364 27344 7392
rect 27338 7352 27344 7364
rect 27396 7352 27402 7404
rect 28000 7401 28028 7500
rect 30006 7420 30012 7472
rect 30064 7420 30070 7472
rect 30116 7460 30144 7500
rect 30282 7488 30288 7540
rect 30340 7528 30346 7540
rect 31297 7531 31355 7537
rect 31297 7528 31309 7531
rect 30340 7500 31309 7528
rect 30340 7488 30346 7500
rect 31297 7497 31309 7500
rect 31343 7497 31355 7531
rect 33686 7528 33692 7540
rect 31297 7491 31355 7497
rect 31404 7500 33692 7528
rect 30374 7460 30380 7472
rect 30116 7432 30380 7460
rect 30374 7420 30380 7432
rect 30432 7460 30438 7472
rect 31404 7460 31432 7500
rect 33686 7488 33692 7500
rect 33744 7488 33750 7540
rect 34330 7488 34336 7540
rect 34388 7528 34394 7540
rect 34517 7531 34575 7537
rect 34517 7528 34529 7531
rect 34388 7500 34529 7528
rect 34388 7488 34394 7500
rect 34517 7497 34529 7500
rect 34563 7497 34575 7531
rect 34517 7491 34575 7497
rect 34790 7460 34796 7472
rect 30432 7432 31432 7460
rect 34270 7432 34796 7460
rect 30432 7420 30438 7432
rect 31404 7401 31432 7432
rect 34790 7420 34796 7432
rect 34848 7420 34854 7472
rect 27985 7395 28043 7401
rect 27985 7361 27997 7395
rect 28031 7361 28043 7395
rect 27985 7355 28043 7361
rect 31389 7395 31447 7401
rect 31389 7361 31401 7395
rect 31435 7361 31447 7395
rect 31389 7355 31447 7361
rect 15286 7324 15292 7336
rect 15199 7296 15292 7324
rect 15286 7284 15292 7296
rect 15344 7324 15350 7336
rect 16022 7324 16028 7336
rect 15344 7296 16028 7324
rect 15344 7284 15350 7296
rect 16022 7284 16028 7296
rect 16080 7284 16086 7336
rect 30466 7324 30472 7336
rect 30427 7296 30472 7324
rect 30466 7284 30472 7296
rect 30524 7284 30530 7336
rect 30745 7327 30803 7333
rect 30745 7293 30757 7327
rect 30791 7324 30803 7327
rect 31846 7324 31852 7336
rect 30791 7296 31852 7324
rect 30791 7293 30803 7296
rect 30745 7287 30803 7293
rect 12158 7188 12164 7200
rect 12119 7160 12164 7188
rect 12158 7148 12164 7160
rect 12216 7148 12222 7200
rect 12802 7148 12808 7200
rect 12860 7188 12866 7200
rect 12897 7191 12955 7197
rect 12897 7188 12909 7191
rect 12860 7160 12909 7188
rect 12860 7148 12866 7160
rect 12897 7157 12909 7160
rect 12943 7157 12955 7191
rect 12897 7151 12955 7157
rect 13541 7191 13599 7197
rect 13541 7157 13553 7191
rect 13587 7188 13599 7191
rect 15470 7188 15476 7200
rect 13587 7160 15476 7188
rect 13587 7157 13599 7160
rect 13541 7151 13599 7157
rect 15470 7148 15476 7160
rect 15528 7148 15534 7200
rect 27154 7188 27160 7200
rect 27115 7160 27160 7188
rect 27154 7148 27160 7160
rect 27212 7148 27218 7200
rect 27890 7188 27896 7200
rect 27851 7160 27896 7188
rect 27890 7148 27896 7160
rect 27948 7148 27954 7200
rect 28994 7188 29000 7200
rect 28955 7160 29000 7188
rect 28994 7148 29000 7160
rect 29052 7148 29058 7200
rect 30282 7148 30288 7200
rect 30340 7188 30346 7200
rect 30760 7188 30788 7287
rect 31846 7284 31852 7296
rect 31904 7284 31910 7336
rect 32674 7284 32680 7336
rect 32732 7324 32738 7336
rect 32769 7327 32827 7333
rect 32769 7324 32781 7327
rect 32732 7296 32781 7324
rect 32732 7284 32738 7296
rect 32769 7293 32781 7296
rect 32815 7293 32827 7327
rect 33042 7324 33048 7336
rect 33003 7296 33048 7324
rect 32769 7287 32827 7293
rect 33042 7284 33048 7296
rect 33100 7284 33106 7336
rect 30340 7160 30788 7188
rect 30340 7148 30346 7160
rect 1104 7098 37628 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 37628 7098
rect 1104 7024 37628 7046
rect 12056 6987 12114 6993
rect 12056 6953 12068 6987
rect 12102 6984 12114 6987
rect 12158 6984 12164 6996
rect 12102 6956 12164 6984
rect 12102 6953 12114 6956
rect 12056 6947 12114 6953
rect 12158 6944 12164 6956
rect 12216 6944 12222 6996
rect 26500 6987 26558 6993
rect 26500 6953 26512 6987
rect 26546 6984 26558 6987
rect 27154 6984 27160 6996
rect 26546 6956 27160 6984
rect 26546 6953 26558 6956
rect 26500 6947 26558 6953
rect 27154 6944 27160 6956
rect 27212 6944 27218 6996
rect 28718 6944 28724 6996
rect 28776 6984 28782 6996
rect 30834 6984 30840 6996
rect 28776 6956 30840 6984
rect 28776 6944 28782 6956
rect 30834 6944 30840 6956
rect 30892 6984 30898 6996
rect 31662 6984 31668 6996
rect 30892 6956 31668 6984
rect 30892 6944 30898 6956
rect 31662 6944 31668 6956
rect 31720 6944 31726 6996
rect 15286 6808 15292 6860
rect 15344 6848 15350 6860
rect 15381 6851 15439 6857
rect 15381 6848 15393 6851
rect 15344 6820 15393 6848
rect 15344 6808 15350 6820
rect 15381 6817 15393 6820
rect 15427 6817 15439 6851
rect 15381 6811 15439 6817
rect 28718 6808 28724 6860
rect 28776 6848 28782 6860
rect 28997 6851 29055 6857
rect 28997 6848 29009 6851
rect 28776 6820 29009 6848
rect 28776 6808 28782 6820
rect 28997 6817 29009 6820
rect 29043 6817 29055 6851
rect 29822 6848 29828 6860
rect 29783 6820 29828 6848
rect 28997 6811 29055 6817
rect 29822 6808 29828 6820
rect 29880 6808 29886 6860
rect 31018 6808 31024 6860
rect 31076 6848 31082 6860
rect 31113 6851 31171 6857
rect 31113 6848 31125 6851
rect 31076 6820 31125 6848
rect 31076 6808 31082 6820
rect 31113 6817 31125 6820
rect 31159 6848 31171 6851
rect 31202 6848 31208 6860
rect 31159 6820 31208 6848
rect 31159 6817 31171 6820
rect 31113 6811 31171 6817
rect 31202 6808 31208 6820
rect 31260 6808 31266 6860
rect 31662 6808 31668 6860
rect 31720 6848 31726 6860
rect 32217 6851 32275 6857
rect 32217 6848 32229 6851
rect 31720 6820 32229 6848
rect 31720 6808 31726 6820
rect 32217 6817 32229 6820
rect 32263 6817 32275 6851
rect 32217 6811 32275 6817
rect 32950 6808 32956 6860
rect 33008 6848 33014 6860
rect 33413 6851 33471 6857
rect 33413 6848 33425 6851
rect 33008 6820 33425 6848
rect 33008 6808 33014 6820
rect 33413 6817 33425 6820
rect 33459 6817 33471 6851
rect 33413 6811 33471 6817
rect 11330 6740 11336 6792
rect 11388 6780 11394 6792
rect 11790 6780 11796 6792
rect 11388 6752 11796 6780
rect 11388 6740 11394 6752
rect 11790 6740 11796 6752
rect 11848 6740 11854 6792
rect 16206 6780 16212 6792
rect 16167 6752 16212 6780
rect 16206 6740 16212 6752
rect 16264 6740 16270 6792
rect 16850 6780 16856 6792
rect 16811 6752 16856 6780
rect 16850 6740 16856 6752
rect 16908 6740 16914 6792
rect 26050 6740 26056 6792
rect 26108 6780 26114 6792
rect 26237 6783 26295 6789
rect 26237 6780 26249 6783
rect 26108 6752 26249 6780
rect 26108 6740 26114 6752
rect 26237 6749 26249 6752
rect 26283 6749 26295 6783
rect 26237 6743 26295 6749
rect 27798 6740 27804 6792
rect 27856 6780 27862 6792
rect 28626 6780 28632 6792
rect 27856 6752 28632 6780
rect 27856 6740 27862 6752
rect 28626 6740 28632 6752
rect 28684 6740 28690 6792
rect 32493 6783 32551 6789
rect 32493 6749 32505 6783
rect 32539 6780 32551 6783
rect 32766 6780 32772 6792
rect 32539 6752 32772 6780
rect 32539 6749 32551 6752
rect 32493 6743 32551 6749
rect 32766 6740 32772 6752
rect 32824 6740 32830 6792
rect 32858 6740 32864 6792
rect 32916 6780 32922 6792
rect 33321 6783 33379 6789
rect 33321 6780 33333 6783
rect 32916 6752 33333 6780
rect 32916 6740 32922 6752
rect 33321 6749 33333 6752
rect 33367 6749 33379 6783
rect 34146 6780 34152 6792
rect 34107 6752 34152 6780
rect 33321 6743 33379 6749
rect 34146 6740 34152 6752
rect 34204 6740 34210 6792
rect 12802 6672 12808 6724
rect 12860 6672 12866 6724
rect 27890 6712 27896 6724
rect 27738 6684 27896 6712
rect 27890 6672 27896 6684
rect 27948 6672 27954 6724
rect 28813 6715 28871 6721
rect 28813 6681 28825 6715
rect 28859 6712 28871 6715
rect 28994 6712 29000 6724
rect 28859 6684 29000 6712
rect 28859 6681 28871 6684
rect 28813 6675 28871 6681
rect 28994 6672 29000 6684
rect 29052 6712 29058 6724
rect 30009 6715 30067 6721
rect 30009 6712 30021 6715
rect 29052 6684 30021 6712
rect 29052 6672 29058 6684
rect 30009 6681 30021 6684
rect 30055 6712 30067 6715
rect 31205 6715 31263 6721
rect 31205 6712 31217 6715
rect 30055 6684 31217 6712
rect 30055 6681 30067 6684
rect 30009 6675 30067 6681
rect 31205 6681 31217 6684
rect 31251 6681 31263 6715
rect 31205 6675 31263 6681
rect 32401 6715 32459 6721
rect 32401 6681 32413 6715
rect 32447 6712 32459 6715
rect 33502 6712 33508 6724
rect 32447 6684 33508 6712
rect 32447 6681 32459 6684
rect 32401 6675 32459 6681
rect 33502 6672 33508 6684
rect 33560 6672 33566 6724
rect 13541 6647 13599 6653
rect 13541 6613 13553 6647
rect 13587 6644 13599 6647
rect 14734 6644 14740 6656
rect 13587 6616 14740 6644
rect 13587 6613 13599 6616
rect 13541 6607 13599 6613
rect 14734 6604 14740 6616
rect 14792 6604 14798 6656
rect 16114 6604 16120 6656
rect 16172 6644 16178 6656
rect 16669 6647 16727 6653
rect 16669 6644 16681 6647
rect 16172 6616 16681 6644
rect 16172 6604 16178 6616
rect 16669 6613 16681 6616
rect 16715 6613 16727 6647
rect 16669 6607 16727 6613
rect 27798 6604 27804 6656
rect 27856 6644 27862 6656
rect 27982 6644 27988 6656
rect 27856 6616 27988 6644
rect 27856 6604 27862 6616
rect 27982 6604 27988 6616
rect 28040 6604 28046 6656
rect 28442 6644 28448 6656
rect 28403 6616 28448 6644
rect 28442 6604 28448 6616
rect 28500 6604 28506 6656
rect 28902 6604 28908 6656
rect 28960 6644 28966 6656
rect 28960 6616 29005 6644
rect 28960 6604 28966 6616
rect 30098 6604 30104 6656
rect 30156 6644 30162 6656
rect 30469 6647 30527 6653
rect 30156 6616 30201 6644
rect 30156 6604 30162 6616
rect 30469 6613 30481 6647
rect 30515 6644 30527 6647
rect 30834 6644 30840 6656
rect 30515 6616 30840 6644
rect 30515 6613 30527 6616
rect 30469 6607 30527 6613
rect 30834 6604 30840 6616
rect 30892 6604 30898 6656
rect 31294 6644 31300 6656
rect 31255 6616 31300 6644
rect 31294 6604 31300 6616
rect 31352 6604 31358 6656
rect 31570 6604 31576 6656
rect 31628 6644 31634 6656
rect 31665 6647 31723 6653
rect 31665 6644 31677 6647
rect 31628 6616 31677 6644
rect 31628 6604 31634 6616
rect 31665 6613 31677 6616
rect 31711 6613 31723 6647
rect 32858 6644 32864 6656
rect 32819 6616 32864 6644
rect 31665 6607 31723 6613
rect 32858 6604 32864 6616
rect 32916 6604 32922 6656
rect 33042 6604 33048 6656
rect 33100 6644 33106 6656
rect 33965 6647 34023 6653
rect 33965 6644 33977 6647
rect 33100 6616 33977 6644
rect 33100 6604 33106 6616
rect 33965 6613 33977 6616
rect 34011 6613 34023 6647
rect 33965 6607 34023 6613
rect 1104 6554 37628 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 35594 6554
rect 35646 6502 35658 6554
rect 35710 6502 35722 6554
rect 35774 6502 35786 6554
rect 35838 6502 35850 6554
rect 35902 6502 37628 6554
rect 1104 6480 37628 6502
rect 12342 6400 12348 6452
rect 12400 6440 12406 6452
rect 12621 6443 12679 6449
rect 12621 6440 12633 6443
rect 12400 6412 12633 6440
rect 12400 6400 12406 6412
rect 12621 6409 12633 6412
rect 12667 6409 12679 6443
rect 12621 6403 12679 6409
rect 13081 6443 13139 6449
rect 13081 6409 13093 6443
rect 13127 6440 13139 6443
rect 14645 6443 14703 6449
rect 14645 6440 14657 6443
rect 13127 6412 14657 6440
rect 13127 6409 13139 6412
rect 13081 6403 13139 6409
rect 14645 6409 14657 6412
rect 14691 6440 14703 6443
rect 14734 6440 14740 6452
rect 14691 6412 14740 6440
rect 14691 6409 14703 6412
rect 14645 6403 14703 6409
rect 14734 6400 14740 6412
rect 14792 6400 14798 6452
rect 16209 6443 16267 6449
rect 16209 6409 16221 6443
rect 16255 6440 16267 6443
rect 16850 6440 16856 6452
rect 16255 6412 16856 6440
rect 16255 6409 16267 6412
rect 16209 6403 16267 6409
rect 16850 6400 16856 6412
rect 16908 6400 16914 6452
rect 27157 6443 27215 6449
rect 27157 6409 27169 6443
rect 27203 6440 27215 6443
rect 27338 6440 27344 6452
rect 27203 6412 27344 6440
rect 27203 6409 27215 6412
rect 27157 6403 27215 6409
rect 27338 6400 27344 6412
rect 27396 6400 27402 6452
rect 27525 6443 27583 6449
rect 27525 6409 27537 6443
rect 27571 6440 27583 6443
rect 28442 6440 28448 6452
rect 27571 6412 28448 6440
rect 27571 6409 27583 6412
rect 27525 6403 27583 6409
rect 28442 6400 28448 6412
rect 28500 6400 28506 6452
rect 28997 6443 29055 6449
rect 28997 6409 29009 6443
rect 29043 6440 29055 6443
rect 29043 6412 30420 6440
rect 29043 6409 29055 6412
rect 28997 6403 29055 6409
rect 15378 6372 15384 6384
rect 14660 6344 15384 6372
rect 11974 6304 11980 6316
rect 11935 6276 11980 6304
rect 11974 6264 11980 6276
rect 12032 6264 12038 6316
rect 12986 6304 12992 6316
rect 12947 6276 12992 6304
rect 12986 6264 12992 6276
rect 13044 6264 13050 6316
rect 13262 6236 13268 6248
rect 13175 6208 13268 6236
rect 13262 6196 13268 6208
rect 13320 6236 13326 6248
rect 14458 6236 14464 6248
rect 13320 6208 14464 6236
rect 13320 6196 13326 6208
rect 14458 6196 14464 6208
rect 14516 6196 14522 6248
rect 14660 6236 14688 6344
rect 15378 6332 15384 6344
rect 15436 6332 15442 6384
rect 17586 6372 17592 6384
rect 16546 6344 17592 6372
rect 14737 6307 14795 6313
rect 14737 6273 14749 6307
rect 14783 6304 14795 6307
rect 15841 6307 15899 6313
rect 15841 6304 15853 6307
rect 14783 6276 15853 6304
rect 14783 6273 14795 6276
rect 14737 6267 14795 6273
rect 15841 6273 15853 6276
rect 15887 6304 15899 6307
rect 16546 6304 16574 6344
rect 17586 6332 17592 6344
rect 17644 6332 17650 6384
rect 29086 6332 29092 6384
rect 29144 6372 29150 6384
rect 30392 6372 30420 6412
rect 30466 6400 30472 6452
rect 30524 6440 30530 6452
rect 31205 6443 31263 6449
rect 31205 6440 31217 6443
rect 30524 6412 31217 6440
rect 30524 6400 30530 6412
rect 31205 6409 31217 6412
rect 31251 6409 31263 6443
rect 31205 6403 31263 6409
rect 31294 6372 31300 6384
rect 29144 6344 29302 6372
rect 30392 6344 31300 6372
rect 29144 6332 29150 6344
rect 31294 6332 31300 6344
rect 31352 6332 31358 6384
rect 33686 6332 33692 6384
rect 33744 6332 33750 6384
rect 15887 6276 16574 6304
rect 16853 6307 16911 6313
rect 15887 6273 15899 6276
rect 15841 6267 15899 6273
rect 16853 6273 16865 6307
rect 16899 6304 16911 6307
rect 17310 6304 17316 6316
rect 16899 6276 17316 6304
rect 16899 6273 16911 6276
rect 16853 6267 16911 6273
rect 17310 6264 17316 6276
rect 17368 6264 17374 6316
rect 26602 6304 26608 6316
rect 26563 6276 26608 6304
rect 26602 6264 26608 6276
rect 26660 6264 26666 6316
rect 28537 6307 28595 6313
rect 28537 6273 28549 6307
rect 28583 6304 28595 6307
rect 29178 6304 29184 6316
rect 28583 6276 29184 6304
rect 28583 6273 28595 6276
rect 28537 6267 28595 6273
rect 29178 6264 29184 6276
rect 29236 6264 29242 6316
rect 30834 6264 30840 6316
rect 30892 6304 30898 6316
rect 31389 6307 31447 6313
rect 31389 6304 31401 6307
rect 30892 6276 31401 6304
rect 30892 6264 30898 6276
rect 31389 6273 31401 6276
rect 31435 6273 31447 6307
rect 31389 6267 31447 6273
rect 34238 6264 34244 6316
rect 34296 6304 34302 6316
rect 35069 6307 35127 6313
rect 35069 6304 35081 6307
rect 34296 6276 35081 6304
rect 34296 6264 34302 6276
rect 35069 6273 35081 6276
rect 35115 6273 35127 6307
rect 35069 6267 35127 6273
rect 14829 6239 14887 6245
rect 14829 6236 14841 6239
rect 14660 6208 14841 6236
rect 14829 6205 14841 6208
rect 14875 6205 14887 6239
rect 14829 6199 14887 6205
rect 13998 6128 14004 6180
rect 14056 6168 14062 6180
rect 14844 6168 14872 6199
rect 15378 6196 15384 6248
rect 15436 6236 15442 6248
rect 15562 6236 15568 6248
rect 15436 6208 15568 6236
rect 15436 6196 15442 6208
rect 15562 6196 15568 6208
rect 15620 6196 15626 6248
rect 15746 6236 15752 6248
rect 15707 6208 15752 6236
rect 15746 6196 15752 6208
rect 15804 6196 15810 6248
rect 27614 6236 27620 6248
rect 27575 6208 27620 6236
rect 27614 6196 27620 6208
rect 27672 6196 27678 6248
rect 27801 6239 27859 6245
rect 27801 6205 27813 6239
rect 27847 6236 27859 6239
rect 29822 6236 29828 6248
rect 27847 6208 29828 6236
rect 27847 6205 27859 6208
rect 27801 6199 27859 6205
rect 29822 6196 29828 6208
rect 29880 6196 29886 6248
rect 30466 6236 30472 6248
rect 30427 6208 30472 6236
rect 30466 6196 30472 6208
rect 30524 6196 30530 6248
rect 30745 6239 30803 6245
rect 30745 6205 30757 6239
rect 30791 6236 30803 6239
rect 32674 6236 32680 6248
rect 30791 6208 32680 6236
rect 30791 6205 30803 6208
rect 30745 6199 30803 6205
rect 14056 6140 14872 6168
rect 14056 6128 14062 6140
rect 11606 6060 11612 6112
rect 11664 6100 11670 6112
rect 11793 6103 11851 6109
rect 11793 6100 11805 6103
rect 11664 6072 11805 6100
rect 11664 6060 11670 6072
rect 11793 6069 11805 6072
rect 11839 6069 11851 6103
rect 11793 6063 11851 6069
rect 14277 6103 14335 6109
rect 14277 6069 14289 6103
rect 14323 6100 14335 6103
rect 14642 6100 14648 6112
rect 14323 6072 14648 6100
rect 14323 6069 14335 6072
rect 14277 6063 14335 6069
rect 14642 6060 14648 6072
rect 14700 6060 14706 6112
rect 16850 6060 16856 6112
rect 16908 6100 16914 6112
rect 16945 6103 17003 6109
rect 16945 6100 16957 6103
rect 16908 6072 16957 6100
rect 16908 6060 16914 6072
rect 16945 6069 16957 6072
rect 16991 6069 17003 6103
rect 16945 6063 17003 6069
rect 26326 6060 26332 6112
rect 26384 6100 26390 6112
rect 26421 6103 26479 6109
rect 26421 6100 26433 6103
rect 26384 6072 26433 6100
rect 26384 6060 26390 6072
rect 26421 6069 26433 6072
rect 26467 6069 26479 6103
rect 28442 6100 28448 6112
rect 28403 6072 28448 6100
rect 26421 6063 26479 6069
rect 28442 6060 28448 6072
rect 28500 6060 28506 6112
rect 30282 6060 30288 6112
rect 30340 6100 30346 6112
rect 30760 6100 30788 6199
rect 32674 6196 32680 6208
rect 32732 6196 32738 6248
rect 32953 6239 33011 6245
rect 32953 6205 32965 6239
rect 32999 6236 33011 6239
rect 32999 6208 34928 6236
rect 32999 6205 33011 6208
rect 32953 6199 33011 6205
rect 34900 6177 34928 6208
rect 34885 6171 34943 6177
rect 34885 6137 34897 6171
rect 34931 6137 34943 6171
rect 34885 6131 34943 6137
rect 30340 6072 30788 6100
rect 30340 6060 30346 6072
rect 33502 6060 33508 6112
rect 33560 6100 33566 6112
rect 34422 6100 34428 6112
rect 33560 6072 34428 6100
rect 33560 6060 33566 6072
rect 34422 6060 34428 6072
rect 34480 6060 34486 6112
rect 1104 6010 37628 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 37628 6010
rect 1104 5936 37628 5958
rect 15013 5899 15071 5905
rect 15013 5865 15025 5899
rect 15059 5896 15071 5899
rect 15930 5896 15936 5908
rect 15059 5868 15936 5896
rect 15059 5865 15071 5868
rect 15013 5859 15071 5865
rect 15930 5856 15936 5868
rect 15988 5856 15994 5908
rect 27706 5856 27712 5908
rect 27764 5896 27770 5908
rect 27801 5899 27859 5905
rect 27801 5896 27813 5899
rect 27764 5868 27813 5896
rect 27764 5856 27770 5868
rect 27801 5865 27813 5868
rect 27847 5896 27859 5899
rect 28902 5896 28908 5908
rect 27847 5868 28908 5896
rect 27847 5865 27859 5868
rect 27801 5859 27859 5865
rect 28902 5856 28908 5868
rect 28960 5856 28966 5908
rect 29086 5896 29092 5908
rect 29047 5868 29092 5896
rect 29086 5856 29092 5868
rect 29144 5856 29150 5908
rect 30006 5856 30012 5908
rect 30064 5896 30070 5908
rect 30101 5899 30159 5905
rect 30101 5896 30113 5899
rect 30064 5868 30113 5896
rect 30064 5856 30070 5868
rect 30101 5865 30113 5868
rect 30147 5865 30159 5899
rect 30101 5859 30159 5865
rect 33873 5899 33931 5905
rect 33873 5865 33885 5899
rect 33919 5896 33931 5899
rect 34238 5896 34244 5908
rect 33919 5868 34244 5896
rect 33919 5865 33931 5868
rect 33873 5859 33931 5865
rect 34238 5856 34244 5868
rect 34296 5856 34302 5908
rect 15470 5828 15476 5840
rect 14568 5800 15476 5828
rect 11606 5760 11612 5772
rect 11567 5732 11612 5760
rect 11606 5720 11612 5732
rect 11664 5720 11670 5772
rect 14458 5760 14464 5772
rect 14419 5732 14464 5760
rect 14458 5720 14464 5732
rect 14516 5720 14522 5772
rect 14568 5769 14596 5800
rect 15470 5788 15476 5800
rect 15528 5828 15534 5840
rect 15746 5828 15752 5840
rect 15528 5800 15752 5828
rect 15528 5788 15534 5800
rect 15746 5788 15752 5800
rect 15804 5788 15810 5840
rect 14553 5763 14611 5769
rect 14553 5729 14565 5763
rect 14599 5729 14611 5763
rect 14553 5723 14611 5729
rect 15286 5720 15292 5772
rect 15344 5760 15350 5772
rect 15562 5760 15568 5772
rect 15344 5732 15568 5760
rect 15344 5720 15350 5732
rect 15562 5720 15568 5732
rect 15620 5760 15626 5772
rect 15841 5763 15899 5769
rect 15841 5760 15853 5763
rect 15620 5732 15853 5760
rect 15620 5720 15626 5732
rect 15841 5729 15853 5732
rect 15887 5729 15899 5763
rect 16114 5760 16120 5772
rect 16075 5732 16120 5760
rect 15841 5723 15899 5729
rect 16114 5720 16120 5732
rect 16172 5720 16178 5772
rect 26326 5760 26332 5772
rect 26287 5732 26332 5760
rect 26326 5720 26332 5732
rect 26384 5720 26390 5772
rect 29730 5720 29736 5772
rect 29788 5760 29794 5772
rect 30282 5760 30288 5772
rect 29788 5732 30288 5760
rect 29788 5720 29794 5732
rect 30282 5720 30288 5732
rect 30340 5760 30346 5772
rect 30929 5763 30987 5769
rect 30929 5760 30941 5763
rect 30340 5732 30941 5760
rect 30340 5720 30346 5732
rect 30929 5729 30941 5732
rect 30975 5729 30987 5763
rect 30929 5723 30987 5729
rect 31202 5720 31208 5772
rect 31260 5760 31266 5772
rect 33229 5763 33287 5769
rect 33229 5760 33241 5763
rect 31260 5732 33241 5760
rect 31260 5720 31266 5732
rect 33229 5729 33241 5732
rect 33275 5729 33287 5763
rect 33229 5723 33287 5729
rect 1765 5695 1823 5701
rect 1765 5661 1777 5695
rect 1811 5692 1823 5695
rect 7006 5692 7012 5704
rect 1811 5664 7012 5692
rect 1811 5661 1823 5664
rect 1765 5655 1823 5661
rect 7006 5652 7012 5664
rect 7064 5652 7070 5704
rect 11330 5692 11336 5704
rect 11291 5664 11336 5692
rect 11330 5652 11336 5664
rect 11388 5652 11394 5704
rect 13541 5695 13599 5701
rect 13541 5661 13553 5695
rect 13587 5692 13599 5695
rect 13722 5692 13728 5704
rect 13587 5664 13728 5692
rect 13587 5661 13599 5664
rect 13541 5655 13599 5661
rect 13722 5652 13728 5664
rect 13780 5652 13786 5704
rect 14642 5692 14648 5704
rect 14603 5664 14648 5692
rect 14642 5652 14648 5664
rect 14700 5652 14706 5704
rect 25038 5652 25044 5704
rect 25096 5692 25102 5704
rect 26050 5692 26056 5704
rect 25096 5664 26056 5692
rect 25096 5652 25102 5664
rect 26050 5652 26056 5664
rect 26108 5652 26114 5704
rect 28442 5692 28448 5704
rect 27462 5664 28448 5692
rect 28442 5652 28448 5664
rect 28500 5652 28506 5704
rect 28997 5695 29055 5701
rect 28997 5661 29009 5695
rect 29043 5692 29055 5695
rect 29178 5692 29184 5704
rect 29043 5664 29184 5692
rect 29043 5661 29055 5664
rect 28997 5655 29055 5661
rect 29178 5652 29184 5664
rect 29236 5652 29242 5704
rect 30009 5695 30067 5701
rect 30009 5661 30021 5695
rect 30055 5692 30067 5695
rect 30374 5692 30380 5704
rect 30055 5664 30380 5692
rect 30055 5661 30067 5664
rect 30009 5655 30067 5661
rect 30374 5652 30380 5664
rect 30432 5652 30438 5704
rect 33502 5692 33508 5704
rect 33463 5664 33508 5692
rect 33502 5652 33508 5664
rect 33560 5652 33566 5704
rect 36906 5692 36912 5704
rect 36867 5664 36912 5692
rect 36906 5652 36912 5664
rect 36964 5652 36970 5704
rect 12618 5584 12624 5636
rect 12676 5584 12682 5636
rect 15286 5624 15292 5636
rect 13740 5596 15292 5624
rect 1578 5556 1584 5568
rect 1539 5528 1584 5556
rect 1578 5516 1584 5528
rect 1636 5516 1642 5568
rect 13078 5556 13084 5568
rect 13039 5528 13084 5556
rect 13078 5516 13084 5528
rect 13136 5516 13142 5568
rect 13740 5565 13768 5596
rect 15286 5584 15292 5596
rect 15344 5584 15350 5636
rect 16850 5584 16856 5636
rect 16908 5584 16914 5636
rect 31202 5624 31208 5636
rect 31163 5596 31208 5624
rect 31202 5584 31208 5596
rect 31260 5584 31266 5636
rect 32582 5624 32588 5636
rect 32430 5596 32588 5624
rect 32582 5584 32588 5596
rect 32640 5584 32646 5636
rect 13725 5559 13783 5565
rect 13725 5525 13737 5559
rect 13771 5525 13783 5559
rect 17586 5556 17592 5568
rect 17547 5528 17592 5556
rect 13725 5519 13783 5525
rect 17586 5516 17592 5528
rect 17644 5516 17650 5568
rect 32677 5559 32735 5565
rect 32677 5525 32689 5559
rect 32723 5556 32735 5559
rect 32766 5556 32772 5568
rect 32723 5528 32772 5556
rect 32723 5525 32735 5528
rect 32677 5519 32735 5525
rect 32766 5516 32772 5528
rect 32824 5556 32830 5568
rect 33413 5559 33471 5565
rect 33413 5556 33425 5559
rect 32824 5528 33425 5556
rect 32824 5516 32830 5528
rect 33413 5525 33425 5528
rect 33459 5525 33471 5559
rect 37090 5556 37096 5568
rect 37051 5528 37096 5556
rect 33413 5519 33471 5525
rect 37090 5516 37096 5528
rect 37148 5516 37154 5568
rect 1104 5466 37628 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 35594 5466
rect 35646 5414 35658 5466
rect 35710 5414 35722 5466
rect 35774 5414 35786 5466
rect 35838 5414 35850 5466
rect 35902 5414 37628 5466
rect 1104 5392 37628 5414
rect 11057 5355 11115 5361
rect 11057 5321 11069 5355
rect 11103 5352 11115 5355
rect 12618 5352 12624 5364
rect 11103 5324 12624 5352
rect 11103 5321 11115 5324
rect 11057 5315 11115 5321
rect 12618 5312 12624 5324
rect 12676 5312 12682 5364
rect 12986 5312 12992 5364
rect 13044 5352 13050 5364
rect 13357 5355 13415 5361
rect 13357 5352 13369 5355
rect 13044 5324 13369 5352
rect 13044 5312 13050 5324
rect 13357 5321 13369 5324
rect 13403 5321 13415 5355
rect 13357 5315 13415 5321
rect 13464 5324 16252 5352
rect 13464 5284 13492 5324
rect 15286 5284 15292 5296
rect 10980 5256 13492 5284
rect 15247 5256 15292 5284
rect 10980 5225 11008 5256
rect 15286 5244 15292 5256
rect 15344 5244 15350 5296
rect 16224 5284 16252 5324
rect 26602 5312 26608 5364
rect 26660 5352 26666 5364
rect 27249 5355 27307 5361
rect 27249 5352 27261 5355
rect 26660 5324 27261 5352
rect 26660 5312 26666 5324
rect 27249 5321 27261 5324
rect 27295 5321 27307 5355
rect 27249 5315 27307 5321
rect 27614 5312 27620 5364
rect 27672 5352 27678 5364
rect 27709 5355 27767 5361
rect 27709 5352 27721 5355
rect 27672 5324 27721 5352
rect 27672 5312 27678 5324
rect 27709 5321 27721 5324
rect 27755 5321 27767 5355
rect 27709 5315 27767 5321
rect 30098 5312 30104 5364
rect 30156 5352 30162 5364
rect 30377 5355 30435 5361
rect 30377 5352 30389 5355
rect 30156 5324 30389 5352
rect 30156 5312 30162 5324
rect 30377 5321 30389 5324
rect 30423 5321 30435 5355
rect 30377 5315 30435 5321
rect 30466 5312 30472 5364
rect 30524 5352 30530 5364
rect 31573 5355 31631 5361
rect 31573 5352 31585 5355
rect 30524 5324 31585 5352
rect 30524 5312 30530 5324
rect 31573 5321 31585 5324
rect 31619 5321 31631 5355
rect 31573 5315 31631 5321
rect 32677 5355 32735 5361
rect 32677 5321 32689 5355
rect 32723 5352 32735 5355
rect 32858 5352 32864 5364
rect 32723 5324 32864 5352
rect 32723 5321 32735 5324
rect 32677 5315 32735 5321
rect 32858 5312 32864 5324
rect 32916 5312 32922 5364
rect 33686 5312 33692 5364
rect 33744 5352 33750 5364
rect 33781 5355 33839 5361
rect 33781 5352 33793 5355
rect 33744 5324 33793 5352
rect 33744 5312 33750 5324
rect 33781 5321 33793 5324
rect 33827 5321 33839 5355
rect 33781 5315 33839 5321
rect 29549 5287 29607 5293
rect 16224 5256 18460 5284
rect 10505 5219 10563 5225
rect 10505 5185 10517 5219
rect 10551 5216 10563 5219
rect 10965 5219 11023 5225
rect 10965 5216 10977 5219
rect 10551 5188 10977 5216
rect 10551 5185 10563 5188
rect 10505 5179 10563 5185
rect 10965 5185 10977 5188
rect 11011 5185 11023 5219
rect 10965 5179 11023 5185
rect 11977 5219 12035 5225
rect 11977 5185 11989 5219
rect 12023 5185 12035 5219
rect 11977 5179 12035 5185
rect 11992 5080 12020 5179
rect 12618 5176 12624 5228
rect 12676 5216 12682 5228
rect 12989 5219 13047 5225
rect 12989 5216 13001 5219
rect 12676 5188 13001 5216
rect 12676 5176 12682 5188
rect 12989 5185 13001 5188
rect 13035 5216 13047 5219
rect 13078 5216 13084 5228
rect 13035 5188 13084 5216
rect 13035 5185 13047 5188
rect 12989 5179 13047 5185
rect 13078 5176 13084 5188
rect 13136 5176 13142 5228
rect 13630 5176 13636 5228
rect 13688 5216 13694 5228
rect 13688 5188 14214 5216
rect 13688 5176 13694 5188
rect 15562 5176 15568 5228
rect 15620 5216 15626 5228
rect 16224 5225 16252 5256
rect 18432 5228 18460 5256
rect 29549 5253 29561 5287
rect 29595 5284 29607 5287
rect 32766 5284 32772 5296
rect 29595 5256 32772 5284
rect 29595 5253 29607 5256
rect 29549 5247 29607 5253
rect 32766 5244 32772 5256
rect 32824 5244 32830 5296
rect 16209 5219 16267 5225
rect 15620 5188 15665 5216
rect 15620 5176 15626 5188
rect 16209 5185 16221 5219
rect 16255 5185 16267 5219
rect 17034 5216 17040 5228
rect 16995 5188 17040 5216
rect 16209 5179 16267 5185
rect 17034 5176 17040 5188
rect 17092 5176 17098 5228
rect 18414 5216 18420 5228
rect 18327 5188 18420 5216
rect 18414 5176 18420 5188
rect 18472 5216 18478 5228
rect 18598 5216 18604 5228
rect 18472 5188 18604 5216
rect 18472 5176 18478 5188
rect 18598 5176 18604 5188
rect 18656 5176 18662 5228
rect 27617 5219 27675 5225
rect 27617 5185 27629 5219
rect 27663 5216 27675 5219
rect 27706 5216 27712 5228
rect 27663 5188 27712 5216
rect 27663 5185 27675 5188
rect 27617 5179 27675 5185
rect 27706 5176 27712 5188
rect 27764 5176 27770 5228
rect 28534 5216 28540 5228
rect 28495 5188 28540 5216
rect 28534 5176 28540 5188
rect 28592 5176 28598 5228
rect 30745 5219 30803 5225
rect 30745 5185 30757 5219
rect 30791 5185 30803 5219
rect 30745 5179 30803 5185
rect 30837 5219 30895 5225
rect 30837 5185 30849 5219
rect 30883 5216 30895 5219
rect 31294 5216 31300 5228
rect 30883 5188 31300 5216
rect 30883 5185 30895 5188
rect 30837 5179 30895 5185
rect 12710 5148 12716 5160
rect 12671 5120 12716 5148
rect 12710 5108 12716 5120
rect 12768 5108 12774 5160
rect 12802 5108 12808 5160
rect 12860 5148 12866 5160
rect 12897 5151 12955 5157
rect 12897 5148 12909 5151
rect 12860 5120 12909 5148
rect 12860 5108 12866 5120
rect 12897 5117 12909 5120
rect 12943 5148 12955 5151
rect 13817 5151 13875 5157
rect 13817 5148 13829 5151
rect 12943 5120 13829 5148
rect 12943 5117 12955 5120
rect 12897 5111 12955 5117
rect 13817 5117 13829 5120
rect 13863 5117 13875 5151
rect 13817 5111 13875 5117
rect 27893 5151 27951 5157
rect 27893 5117 27905 5151
rect 27939 5117 27951 5151
rect 29638 5148 29644 5160
rect 29599 5120 29644 5148
rect 27893 5111 27951 5117
rect 13538 5080 13544 5092
rect 11992 5052 13544 5080
rect 13538 5040 13544 5052
rect 13596 5040 13602 5092
rect 27908 5080 27936 5111
rect 29638 5108 29644 5120
rect 29696 5108 29702 5160
rect 29825 5151 29883 5157
rect 29825 5117 29837 5151
rect 29871 5148 29883 5151
rect 29871 5120 30604 5148
rect 29871 5117 29883 5120
rect 29825 5111 29883 5117
rect 28810 5080 28816 5092
rect 27908 5052 28816 5080
rect 28810 5040 28816 5052
rect 28868 5080 28874 5092
rect 30006 5080 30012 5092
rect 28868 5052 30012 5080
rect 28868 5040 28874 5052
rect 30006 5040 30012 5052
rect 30064 5040 30070 5092
rect 10413 5015 10471 5021
rect 10413 4981 10425 5015
rect 10459 5012 10471 5015
rect 10870 5012 10876 5024
rect 10459 4984 10876 5012
rect 10459 4981 10471 4984
rect 10413 4975 10471 4981
rect 10870 4972 10876 4984
rect 10928 4972 10934 5024
rect 12066 5012 12072 5024
rect 12027 4984 12072 5012
rect 12066 4972 12072 4984
rect 12124 4972 12130 5024
rect 15470 4972 15476 5024
rect 15528 5012 15534 5024
rect 16117 5015 16175 5021
rect 16117 5012 16129 5015
rect 15528 4984 16129 5012
rect 15528 4972 15534 4984
rect 16117 4981 16129 4984
rect 16163 4981 16175 5015
rect 16850 5012 16856 5024
rect 16811 4984 16856 5012
rect 16117 4975 16175 4981
rect 16850 4972 16856 4984
rect 16908 4972 16914 5024
rect 18138 4972 18144 5024
rect 18196 5012 18202 5024
rect 18325 5015 18383 5021
rect 18325 5012 18337 5015
rect 18196 4984 18337 5012
rect 18196 4972 18202 4984
rect 18325 4981 18337 4984
rect 18371 4981 18383 5015
rect 18325 4975 18383 4981
rect 28721 5015 28779 5021
rect 28721 4981 28733 5015
rect 28767 5012 28779 5015
rect 28994 5012 29000 5024
rect 28767 4984 29000 5012
rect 28767 4981 28779 4984
rect 28721 4975 28779 4981
rect 28994 4972 29000 4984
rect 29052 4972 29058 5024
rect 29178 5012 29184 5024
rect 29139 4984 29184 5012
rect 29178 4972 29184 4984
rect 29236 4972 29242 5024
rect 30576 5012 30604 5120
rect 30760 5080 30788 5179
rect 31294 5176 31300 5188
rect 31352 5176 31358 5228
rect 31570 5176 31576 5228
rect 31628 5216 31634 5228
rect 31757 5219 31815 5225
rect 31757 5216 31769 5219
rect 31628 5188 31769 5216
rect 31628 5176 31634 5188
rect 31757 5185 31769 5188
rect 31803 5185 31815 5219
rect 31757 5179 31815 5185
rect 33689 5219 33747 5225
rect 33689 5185 33701 5219
rect 33735 5216 33747 5219
rect 33778 5216 33784 5228
rect 33735 5188 33784 5216
rect 33735 5185 33747 5188
rect 33689 5179 33747 5185
rect 33778 5176 33784 5188
rect 33836 5176 33842 5228
rect 30926 5148 30932 5160
rect 30887 5120 30932 5148
rect 30926 5108 30932 5120
rect 30984 5148 30990 5160
rect 31662 5148 31668 5160
rect 30984 5120 31668 5148
rect 30984 5108 30990 5120
rect 31662 5108 31668 5120
rect 31720 5108 31726 5160
rect 32490 5108 32496 5160
rect 32548 5148 32554 5160
rect 32858 5148 32864 5160
rect 32548 5120 32864 5148
rect 32548 5108 32554 5120
rect 32858 5108 32864 5120
rect 32916 5108 32922 5160
rect 34790 5080 34796 5092
rect 30760 5052 34796 5080
rect 34790 5040 34796 5052
rect 34848 5040 34854 5092
rect 30926 5012 30932 5024
rect 30576 4984 30932 5012
rect 30926 4972 30932 4984
rect 30984 4972 30990 5024
rect 32122 4972 32128 5024
rect 32180 5012 32186 5024
rect 32309 5015 32367 5021
rect 32309 5012 32321 5015
rect 32180 4984 32321 5012
rect 32180 4972 32186 4984
rect 32309 4981 32321 4984
rect 32355 4981 32367 5015
rect 32309 4975 32367 4981
rect 1104 4922 37628 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 37628 4922
rect 1104 4848 37628 4870
rect 11974 4768 11980 4820
rect 12032 4808 12038 4820
rect 12161 4811 12219 4817
rect 12161 4808 12173 4811
rect 12032 4780 12173 4808
rect 12032 4768 12038 4780
rect 12161 4777 12173 4780
rect 12207 4777 12219 4811
rect 13630 4808 13636 4820
rect 13591 4780 13636 4808
rect 12161 4771 12219 4777
rect 13630 4768 13636 4780
rect 13688 4768 13694 4820
rect 13722 4768 13728 4820
rect 13780 4808 13786 4820
rect 14277 4811 14335 4817
rect 14277 4808 14289 4811
rect 13780 4780 14289 4808
rect 13780 4768 13786 4780
rect 14277 4777 14289 4780
rect 14323 4777 14335 4811
rect 18690 4808 18696 4820
rect 18603 4780 18696 4808
rect 14277 4771 14335 4777
rect 10965 4743 11023 4749
rect 10965 4709 10977 4743
rect 11011 4709 11023 4743
rect 18616 4740 18644 4780
rect 18690 4768 18696 4780
rect 18748 4808 18754 4820
rect 18748 4780 22692 4808
rect 18748 4768 18754 4780
rect 10965 4703 11023 4709
rect 17328 4712 18644 4740
rect 10321 4607 10379 4613
rect 10321 4573 10333 4607
rect 10367 4604 10379 4607
rect 10980 4604 11008 4703
rect 11609 4675 11667 4681
rect 11609 4641 11621 4675
rect 11655 4672 11667 4675
rect 12805 4675 12863 4681
rect 12805 4672 12817 4675
rect 11655 4644 12817 4672
rect 11655 4641 11667 4644
rect 11609 4635 11667 4641
rect 12805 4641 12817 4644
rect 12851 4672 12863 4675
rect 13262 4672 13268 4684
rect 12851 4644 13268 4672
rect 12851 4641 12863 4644
rect 12805 4635 12863 4641
rect 13262 4632 13268 4644
rect 13320 4632 13326 4684
rect 14734 4672 14740 4684
rect 14695 4644 14740 4672
rect 14734 4632 14740 4644
rect 14792 4632 14798 4684
rect 14826 4632 14832 4684
rect 14884 4672 14890 4684
rect 15378 4672 15384 4684
rect 14884 4644 15384 4672
rect 14884 4632 14890 4644
rect 15378 4632 15384 4644
rect 15436 4632 15442 4684
rect 16485 4675 16543 4681
rect 16485 4641 16497 4675
rect 16531 4672 16543 4675
rect 17328 4672 17356 4712
rect 16531 4644 17356 4672
rect 16531 4641 16543 4644
rect 16485 4635 16543 4641
rect 17402 4632 17408 4684
rect 17460 4632 17466 4684
rect 18616 4681 18644 4712
rect 22465 4743 22523 4749
rect 22465 4709 22477 4743
rect 22511 4709 22523 4743
rect 22465 4703 22523 4709
rect 18601 4675 18659 4681
rect 18601 4641 18613 4675
rect 18647 4641 18659 4675
rect 22370 4672 22376 4684
rect 18601 4635 18659 4641
rect 19812 4644 22376 4672
rect 13538 4604 13544 4616
rect 10367 4576 11008 4604
rect 13499 4576 13544 4604
rect 10367 4573 10379 4576
rect 10321 4567 10379 4573
rect 13538 4564 13544 4576
rect 13596 4564 13602 4616
rect 17129 4607 17187 4613
rect 17129 4573 17141 4607
rect 17175 4604 17187 4607
rect 17420 4604 17448 4632
rect 19812 4604 19840 4644
rect 22370 4632 22376 4644
rect 22428 4632 22434 4684
rect 19978 4604 19984 4616
rect 17175 4576 19840 4604
rect 19939 4576 19984 4604
rect 17175 4573 17187 4576
rect 17129 4567 17187 4573
rect 19978 4564 19984 4576
rect 20036 4564 20042 4616
rect 20625 4607 20683 4613
rect 20625 4573 20637 4607
rect 20671 4573 20683 4607
rect 20625 4567 20683 4573
rect 21821 4607 21879 4613
rect 21821 4573 21833 4607
rect 21867 4604 21879 4607
rect 22480 4604 22508 4703
rect 22664 4684 22692 4780
rect 28736 4780 31156 4808
rect 22646 4632 22652 4684
rect 22704 4672 22710 4684
rect 28736 4681 28764 4780
rect 23109 4675 23167 4681
rect 23109 4672 23121 4675
rect 22704 4644 23121 4672
rect 22704 4632 22710 4644
rect 23109 4641 23121 4644
rect 23155 4672 23167 4675
rect 28721 4675 28779 4681
rect 28721 4672 28733 4675
rect 23155 4644 28733 4672
rect 23155 4641 23167 4644
rect 23109 4635 23167 4641
rect 28721 4641 28733 4644
rect 28767 4641 28779 4675
rect 28721 4635 28779 4641
rect 28994 4632 29000 4684
rect 29052 4672 29058 4684
rect 30009 4675 30067 4681
rect 30009 4672 30021 4675
rect 29052 4644 30021 4672
rect 29052 4632 29058 4644
rect 30009 4641 30021 4644
rect 30055 4641 30067 4675
rect 31128 4672 31156 4780
rect 31202 4768 31208 4820
rect 31260 4808 31266 4820
rect 31941 4811 31999 4817
rect 31941 4808 31953 4811
rect 31260 4780 31953 4808
rect 31260 4768 31266 4780
rect 31941 4777 31953 4780
rect 31987 4777 31999 4811
rect 31941 4771 31999 4777
rect 32582 4768 32588 4820
rect 32640 4808 32646 4820
rect 32677 4811 32735 4817
rect 32677 4808 32689 4811
rect 32640 4780 32689 4808
rect 32640 4768 32646 4780
rect 32677 4777 32689 4780
rect 32723 4777 32735 4811
rect 32677 4771 32735 4777
rect 31478 4740 31484 4752
rect 31391 4712 31484 4740
rect 31478 4700 31484 4712
rect 31536 4740 31542 4752
rect 36906 4740 36912 4752
rect 31536 4712 36912 4740
rect 31536 4700 31542 4712
rect 36906 4700 36912 4712
rect 36964 4700 36970 4752
rect 32858 4672 32864 4684
rect 31128 4644 32864 4672
rect 30009 4635 30067 4641
rect 32858 4632 32864 4644
rect 32916 4632 32922 4684
rect 23842 4604 23848 4616
rect 21867 4576 22508 4604
rect 22572 4576 23848 4604
rect 21867 4573 21879 4576
rect 21821 4567 21879 4573
rect 11333 4539 11391 4545
rect 11333 4505 11345 4539
rect 11379 4536 11391 4539
rect 12894 4536 12900 4548
rect 11379 4508 12900 4536
rect 11379 4505 11391 4508
rect 11333 4499 11391 4505
rect 12894 4496 12900 4508
rect 12952 4496 12958 4548
rect 14550 4496 14556 4548
rect 14608 4536 14614 4548
rect 16393 4539 16451 4545
rect 16393 4536 16405 4539
rect 14608 4508 16405 4536
rect 14608 4496 14614 4508
rect 16393 4505 16405 4508
rect 16439 4505 16451 4539
rect 16393 4499 16451 4505
rect 17310 4496 17316 4548
rect 17368 4536 17374 4548
rect 17405 4539 17463 4545
rect 17405 4536 17417 4539
rect 17368 4508 17417 4536
rect 17368 4496 17374 4508
rect 17405 4505 17417 4508
rect 17451 4505 17463 4539
rect 17405 4499 17463 4505
rect 17954 4496 17960 4548
rect 18012 4536 18018 4548
rect 18012 4508 18552 4536
rect 18012 4496 18018 4508
rect 10505 4471 10563 4477
rect 10505 4437 10517 4471
rect 10551 4468 10563 4471
rect 10778 4468 10784 4480
rect 10551 4440 10784 4468
rect 10551 4437 10563 4440
rect 10505 4431 10563 4437
rect 10778 4428 10784 4440
rect 10836 4428 10842 4480
rect 11425 4471 11483 4477
rect 11425 4437 11437 4471
rect 11471 4468 11483 4471
rect 12342 4468 12348 4480
rect 11471 4440 12348 4468
rect 11471 4437 11483 4440
rect 11425 4431 11483 4437
rect 12342 4428 12348 4440
rect 12400 4428 12406 4480
rect 12526 4468 12532 4480
rect 12487 4440 12532 4468
rect 12526 4428 12532 4440
rect 12584 4428 12590 4480
rect 12618 4428 12624 4480
rect 12676 4468 12682 4480
rect 12676 4440 12721 4468
rect 12676 4428 12682 4440
rect 12802 4428 12808 4480
rect 12860 4468 12866 4480
rect 14645 4471 14703 4477
rect 14645 4468 14657 4471
rect 12860 4440 14657 4468
rect 12860 4428 12866 4440
rect 14645 4437 14657 4440
rect 14691 4437 14703 4471
rect 15930 4468 15936 4480
rect 15891 4440 15936 4468
rect 14645 4431 14703 4437
rect 15930 4428 15936 4440
rect 15988 4428 15994 4480
rect 16206 4428 16212 4480
rect 16264 4468 16270 4480
rect 16301 4471 16359 4477
rect 16301 4468 16313 4471
rect 16264 4440 16313 4468
rect 16264 4428 16270 4440
rect 16301 4437 16313 4440
rect 16347 4437 16359 4471
rect 18046 4468 18052 4480
rect 18007 4440 18052 4468
rect 16301 4431 16359 4437
rect 18046 4428 18052 4440
rect 18104 4428 18110 4480
rect 18414 4468 18420 4480
rect 18375 4440 18420 4468
rect 18414 4428 18420 4440
rect 18472 4428 18478 4480
rect 18524 4477 18552 4508
rect 18598 4496 18604 4548
rect 18656 4536 18662 4548
rect 20640 4536 20668 4567
rect 22572 4536 22600 4576
rect 23842 4564 23848 4576
rect 23900 4564 23906 4616
rect 27709 4607 27767 4613
rect 27709 4573 27721 4607
rect 27755 4604 27767 4607
rect 28537 4607 28595 4613
rect 27755 4576 28212 4604
rect 27755 4573 27767 4576
rect 27709 4567 27767 4573
rect 18656 4508 22600 4536
rect 22833 4539 22891 4545
rect 18656 4496 18662 4508
rect 22833 4505 22845 4539
rect 22879 4536 22891 4539
rect 23290 4536 23296 4548
rect 22879 4508 23296 4536
rect 22879 4505 22891 4508
rect 22833 4499 22891 4505
rect 23290 4496 23296 4508
rect 23348 4496 23354 4548
rect 18509 4471 18567 4477
rect 18509 4437 18521 4471
rect 18555 4468 18567 4471
rect 18874 4468 18880 4480
rect 18555 4440 18880 4468
rect 18555 4437 18567 4440
rect 18509 4431 18567 4437
rect 18874 4428 18880 4440
rect 18932 4428 18938 4480
rect 19610 4428 19616 4480
rect 19668 4468 19674 4480
rect 19797 4471 19855 4477
rect 19797 4468 19809 4471
rect 19668 4440 19809 4468
rect 19668 4428 19674 4440
rect 19797 4437 19809 4440
rect 19843 4437 19855 4471
rect 19797 4431 19855 4437
rect 20533 4471 20591 4477
rect 20533 4437 20545 4471
rect 20579 4468 20591 4471
rect 20622 4468 20628 4480
rect 20579 4440 20628 4468
rect 20579 4437 20591 4440
rect 20533 4431 20591 4437
rect 20622 4428 20628 4440
rect 20680 4428 20686 4480
rect 22002 4468 22008 4480
rect 21963 4440 22008 4468
rect 22002 4428 22008 4440
rect 22060 4428 22066 4480
rect 22922 4468 22928 4480
rect 22883 4440 22928 4468
rect 22922 4428 22928 4440
rect 22980 4428 22986 4480
rect 27522 4468 27528 4480
rect 27483 4440 27528 4468
rect 27522 4428 27528 4440
rect 27580 4428 27586 4480
rect 28184 4477 28212 4576
rect 28537 4573 28549 4607
rect 28583 4604 28595 4607
rect 29178 4604 29184 4616
rect 28583 4576 29184 4604
rect 28583 4573 28595 4576
rect 28537 4567 28595 4573
rect 29178 4564 29184 4576
rect 29236 4564 29242 4616
rect 29730 4604 29736 4616
rect 29691 4576 29736 4604
rect 29730 4564 29736 4576
rect 29788 4564 29794 4616
rect 32122 4604 32128 4616
rect 32083 4576 32128 4604
rect 32122 4564 32128 4576
rect 32180 4564 32186 4616
rect 32766 4604 32772 4616
rect 32727 4576 32772 4604
rect 32766 4564 32772 4576
rect 32824 4604 32830 4616
rect 32950 4604 32956 4616
rect 32824 4576 32956 4604
rect 32824 4564 32830 4576
rect 32950 4564 32956 4576
rect 33008 4564 33014 4616
rect 30742 4496 30748 4548
rect 30800 4496 30806 4548
rect 28169 4471 28227 4477
rect 28169 4437 28181 4471
rect 28215 4437 28227 4471
rect 28169 4431 28227 4437
rect 28442 4428 28448 4480
rect 28500 4468 28506 4480
rect 28629 4471 28687 4477
rect 28629 4468 28641 4471
rect 28500 4440 28641 4468
rect 28500 4428 28506 4440
rect 28629 4437 28641 4440
rect 28675 4437 28687 4471
rect 28629 4431 28687 4437
rect 1104 4378 37628 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 35594 4378
rect 35646 4326 35658 4378
rect 35710 4326 35722 4378
rect 35774 4326 35786 4378
rect 35838 4326 35850 4378
rect 35902 4326 37628 4378
rect 1104 4304 37628 4326
rect 12437 4267 12495 4273
rect 12437 4264 12449 4267
rect 12268 4236 12449 4264
rect 10781 4199 10839 4205
rect 10781 4165 10793 4199
rect 10827 4165 10839 4199
rect 10781 4159 10839 4165
rect 10796 4128 10824 4159
rect 10962 4128 10968 4140
rect 10796 4100 10968 4128
rect 10962 4088 10968 4100
rect 11020 4128 11026 4140
rect 12268 4128 12296 4236
rect 12437 4233 12449 4236
rect 12483 4233 12495 4267
rect 12437 4227 12495 4233
rect 12526 4224 12532 4276
rect 12584 4264 12590 4276
rect 12897 4267 12955 4273
rect 12897 4264 12909 4267
rect 12584 4236 12909 4264
rect 12584 4224 12590 4236
rect 12897 4233 12909 4236
rect 12943 4233 12955 4267
rect 12897 4227 12955 4233
rect 15654 4224 15660 4276
rect 15712 4224 15718 4276
rect 18874 4264 18880 4276
rect 18835 4236 18880 4264
rect 18874 4224 18880 4236
rect 18932 4224 18938 4276
rect 23106 4224 23112 4276
rect 23164 4264 23170 4276
rect 24581 4267 24639 4273
rect 23164 4236 23612 4264
rect 23164 4224 23170 4236
rect 13725 4199 13783 4205
rect 11020 4100 12296 4128
rect 12360 4168 12756 4196
rect 11020 4088 11026 4100
rect 12360 4069 12388 4168
rect 12728 4140 12756 4168
rect 13725 4165 13737 4199
rect 13771 4196 13783 4199
rect 14550 4196 14556 4208
rect 13771 4168 14556 4196
rect 13771 4165 13783 4168
rect 13725 4159 13783 4165
rect 14550 4156 14556 4168
rect 14608 4156 14614 4208
rect 15470 4156 15476 4208
rect 15528 4156 15534 4208
rect 15672 4196 15700 4224
rect 15672 4168 16344 4196
rect 16316 4140 16344 4168
rect 18138 4156 18144 4208
rect 18196 4156 18202 4208
rect 19610 4196 19616 4208
rect 19571 4168 19616 4196
rect 19610 4156 19616 4168
rect 19668 4156 19674 4208
rect 20622 4156 20628 4208
rect 20680 4156 20686 4208
rect 22002 4156 22008 4208
rect 22060 4196 22066 4208
rect 22281 4199 22339 4205
rect 22281 4196 22293 4199
rect 22060 4168 22293 4196
rect 22060 4156 22066 4168
rect 22281 4165 22293 4168
rect 22327 4165 22339 4199
rect 22281 4159 22339 4165
rect 12434 4088 12440 4140
rect 12492 4128 12498 4140
rect 12529 4131 12587 4137
rect 12529 4128 12541 4131
rect 12492 4100 12541 4128
rect 12492 4088 12498 4100
rect 12529 4097 12541 4100
rect 12575 4097 12587 4131
rect 12529 4091 12587 4097
rect 12710 4088 12716 4140
rect 12768 4128 12774 4140
rect 12768 4100 14044 4128
rect 12768 4088 12774 4100
rect 14016 4072 14044 4100
rect 16298 4088 16304 4140
rect 16356 4128 16362 4140
rect 16356 4100 16574 4128
rect 16356 4088 16362 4100
rect 10873 4063 10931 4069
rect 10873 4029 10885 4063
rect 10919 4029 10931 4063
rect 10873 4023 10931 4029
rect 11057 4063 11115 4069
rect 11057 4029 11069 4063
rect 11103 4029 11115 4063
rect 11057 4023 11115 4029
rect 12345 4063 12403 4069
rect 12345 4029 12357 4063
rect 12391 4029 12403 4063
rect 13262 4060 13268 4072
rect 12345 4023 12403 4029
rect 12820 4032 13268 4060
rect 9858 3884 9864 3936
rect 9916 3924 9922 3936
rect 10413 3927 10471 3933
rect 10413 3924 10425 3927
rect 9916 3896 10425 3924
rect 9916 3884 9922 3896
rect 10413 3893 10425 3896
rect 10459 3893 10471 3927
rect 10888 3924 10916 4023
rect 11072 3992 11100 4023
rect 12820 3992 12848 4032
rect 13262 4020 13268 4032
rect 13320 4020 13326 4072
rect 13817 4063 13875 4069
rect 13817 4029 13829 4063
rect 13863 4029 13875 4063
rect 13998 4060 14004 4072
rect 13959 4032 14004 4060
rect 13817 4023 13875 4029
rect 11072 3964 12848 3992
rect 12894 3952 12900 4004
rect 12952 3992 12958 4004
rect 13357 3995 13415 4001
rect 13357 3992 13369 3995
rect 12952 3964 13369 3992
rect 12952 3952 12958 3964
rect 13357 3961 13369 3964
rect 13403 3961 13415 3995
rect 13357 3955 13415 3961
rect 12618 3924 12624 3936
rect 10888 3896 12624 3924
rect 10413 3887 10471 3893
rect 12618 3884 12624 3896
rect 12676 3884 12682 3936
rect 12986 3884 12992 3936
rect 13044 3924 13050 3936
rect 13832 3924 13860 4023
rect 13998 4020 14004 4032
rect 14056 4020 14062 4072
rect 14550 4060 14556 4072
rect 14511 4032 14556 4060
rect 14550 4020 14556 4032
rect 14608 4020 14614 4072
rect 16022 4060 16028 4072
rect 15983 4032 16028 4060
rect 16022 4020 16028 4032
rect 16080 4020 16086 4072
rect 16546 4060 16574 4100
rect 23382 4088 23388 4140
rect 23440 4088 23446 4140
rect 23584 4128 23612 4236
rect 24581 4233 24593 4267
rect 24627 4264 24639 4267
rect 28442 4264 28448 4276
rect 24627 4236 28448 4264
rect 24627 4233 24639 4236
rect 24581 4227 24639 4233
rect 28442 4224 28448 4236
rect 28500 4224 28506 4276
rect 28534 4224 28540 4276
rect 28592 4264 28598 4276
rect 29457 4267 29515 4273
rect 29457 4264 29469 4267
rect 28592 4236 29469 4264
rect 28592 4224 28598 4236
rect 29457 4233 29469 4236
rect 29503 4233 29515 4267
rect 29457 4227 29515 4233
rect 29638 4224 29644 4276
rect 29696 4264 29702 4276
rect 29825 4267 29883 4273
rect 29825 4264 29837 4267
rect 29696 4236 29837 4264
rect 29696 4224 29702 4236
rect 29825 4233 29837 4236
rect 29871 4264 29883 4267
rect 31478 4264 31484 4276
rect 29871 4236 31484 4264
rect 29871 4233 29883 4236
rect 29825 4227 29883 4233
rect 31478 4224 31484 4236
rect 31536 4224 31542 4276
rect 27522 4196 27528 4208
rect 27483 4168 27528 4196
rect 27522 4156 27528 4168
rect 27580 4156 27586 4208
rect 28074 4156 28080 4208
rect 28132 4156 28138 4208
rect 23584 4100 24808 4128
rect 17129 4063 17187 4069
rect 17129 4060 17141 4063
rect 16546 4032 17141 4060
rect 17129 4029 17141 4032
rect 17175 4029 17187 4063
rect 17129 4023 17187 4029
rect 17405 4063 17463 4069
rect 17405 4029 17417 4063
rect 17451 4060 17463 4063
rect 17494 4060 17500 4072
rect 17451 4032 17500 4060
rect 17451 4029 17463 4032
rect 17405 4023 17463 4029
rect 13044 3896 13860 3924
rect 17144 3924 17172 4023
rect 17494 4020 17500 4032
rect 17552 4020 17558 4072
rect 19337 4063 19395 4069
rect 19337 4029 19349 4063
rect 19383 4029 19395 4063
rect 22002 4060 22008 4072
rect 21963 4032 22008 4060
rect 19337 4023 19395 4029
rect 19352 3992 19380 4023
rect 22002 4020 22008 4032
rect 22060 4020 22066 4072
rect 22922 4020 22928 4072
rect 22980 4060 22986 4072
rect 24780 4069 24808 4100
rect 28902 4088 28908 4140
rect 28960 4128 28966 4140
rect 30653 4131 30711 4137
rect 30653 4128 30665 4131
rect 28960 4100 30665 4128
rect 28960 4088 28966 4100
rect 30653 4097 30665 4100
rect 30699 4097 30711 4131
rect 30653 4091 30711 4097
rect 23753 4063 23811 4069
rect 23753 4060 23765 4063
rect 22980 4032 23765 4060
rect 22980 4020 22986 4032
rect 23753 4029 23765 4032
rect 23799 4029 23811 4063
rect 23753 4023 23811 4029
rect 24673 4063 24731 4069
rect 24673 4029 24685 4063
rect 24719 4029 24731 4063
rect 24673 4023 24731 4029
rect 24765 4063 24823 4069
rect 24765 4029 24777 4063
rect 24811 4029 24823 4063
rect 24765 4023 24823 4029
rect 27249 4063 27307 4069
rect 27249 4029 27261 4063
rect 27295 4029 27307 4063
rect 27249 4023 27307 4029
rect 18432 3964 19380 3992
rect 18432 3924 18460 3964
rect 23290 3952 23296 4004
rect 23348 3992 23354 4004
rect 24213 3995 24271 4001
rect 24213 3992 24225 3995
rect 23348 3964 24225 3992
rect 23348 3952 23354 3964
rect 24213 3961 24225 3964
rect 24259 3961 24271 3995
rect 24213 3955 24271 3961
rect 17144 3896 18460 3924
rect 13044 3884 13050 3896
rect 20622 3884 20628 3936
rect 20680 3924 20686 3936
rect 21085 3927 21143 3933
rect 21085 3924 21097 3927
rect 20680 3896 21097 3924
rect 20680 3884 20686 3896
rect 21085 3893 21097 3896
rect 21131 3893 21143 3927
rect 21085 3887 21143 3893
rect 23014 3884 23020 3936
rect 23072 3924 23078 3936
rect 24688 3924 24716 4023
rect 27154 3924 27160 3936
rect 23072 3896 27160 3924
rect 23072 3884 23078 3896
rect 27154 3884 27160 3896
rect 27212 3884 27218 3936
rect 27264 3924 27292 4023
rect 28534 4020 28540 4072
rect 28592 4060 28598 4072
rect 28997 4063 29055 4069
rect 28997 4060 29009 4063
rect 28592 4032 29009 4060
rect 28592 4020 28598 4032
rect 28997 4029 29009 4032
rect 29043 4060 29055 4063
rect 29917 4063 29975 4069
rect 29917 4060 29929 4063
rect 29043 4032 29929 4060
rect 29043 4029 29055 4032
rect 28997 4023 29055 4029
rect 29917 4029 29929 4032
rect 29963 4029 29975 4063
rect 29917 4023 29975 4029
rect 30006 4020 30012 4072
rect 30064 4060 30070 4072
rect 30668 4060 30696 4091
rect 30742 4088 30748 4140
rect 30800 4128 30806 4140
rect 30800 4100 30845 4128
rect 30800 4088 30806 4100
rect 33778 4060 33784 4072
rect 30064 4032 30109 4060
rect 30668 4032 33784 4060
rect 30064 4020 30070 4032
rect 33778 4020 33784 4032
rect 33836 4020 33842 4072
rect 29730 3992 29736 4004
rect 28920 3964 29736 3992
rect 28920 3924 28948 3964
rect 29730 3952 29736 3964
rect 29788 3952 29794 4004
rect 27264 3896 28948 3924
rect 1104 3834 37628 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 37628 3834
rect 1104 3760 37628 3782
rect 12253 3723 12311 3729
rect 12253 3689 12265 3723
rect 12299 3720 12311 3723
rect 12342 3720 12348 3732
rect 12299 3692 12348 3720
rect 12299 3689 12311 3692
rect 12253 3683 12311 3689
rect 12342 3680 12348 3692
rect 12400 3720 12406 3732
rect 12400 3692 13308 3720
rect 12400 3680 12406 3692
rect 11882 3612 11888 3664
rect 11940 3652 11946 3664
rect 12986 3652 12992 3664
rect 11940 3624 12992 3652
rect 11940 3612 11946 3624
rect 12986 3612 12992 3624
rect 13044 3612 13050 3664
rect 10505 3587 10563 3593
rect 10505 3553 10517 3587
rect 10551 3584 10563 3587
rect 11330 3584 11336 3596
rect 10551 3556 11336 3584
rect 10551 3553 10563 3556
rect 10505 3547 10563 3553
rect 11330 3544 11336 3556
rect 11388 3584 11394 3596
rect 12158 3584 12164 3596
rect 11388 3556 12164 3584
rect 11388 3544 11394 3556
rect 12158 3544 12164 3556
rect 12216 3544 12222 3596
rect 9858 3516 9864 3528
rect 9819 3488 9864 3516
rect 9858 3476 9864 3488
rect 9916 3476 9922 3528
rect 12066 3476 12072 3528
rect 12124 3516 12130 3528
rect 13078 3516 13084 3528
rect 12124 3488 13084 3516
rect 12124 3476 12130 3488
rect 13078 3476 13084 3488
rect 13136 3476 13142 3528
rect 10778 3448 10784 3460
rect 10739 3420 10784 3448
rect 10778 3408 10784 3420
rect 10836 3408 10842 3460
rect 10870 3408 10876 3460
rect 10928 3448 10934 3460
rect 12894 3448 12900 3460
rect 10928 3420 11270 3448
rect 12268 3420 12900 3448
rect 10928 3408 10934 3420
rect 10045 3383 10103 3389
rect 10045 3349 10057 3383
rect 10091 3380 10103 3383
rect 12268 3380 12296 3420
rect 12894 3408 12900 3420
rect 12952 3408 12958 3460
rect 10091 3352 12296 3380
rect 10091 3349 10103 3352
rect 10045 3343 10103 3349
rect 12342 3340 12348 3392
rect 12400 3380 12406 3392
rect 12713 3383 12771 3389
rect 12713 3380 12725 3383
rect 12400 3352 12725 3380
rect 12400 3340 12406 3352
rect 12713 3349 12725 3352
rect 12759 3349 12771 3383
rect 12713 3343 12771 3349
rect 12986 3340 12992 3392
rect 13044 3380 13050 3392
rect 13081 3383 13139 3389
rect 13081 3380 13093 3383
rect 13044 3352 13093 3380
rect 13044 3340 13050 3352
rect 13081 3349 13093 3352
rect 13127 3349 13139 3383
rect 13081 3343 13139 3349
rect 13173 3383 13231 3389
rect 13173 3349 13185 3383
rect 13219 3380 13231 3383
rect 13280 3380 13308 3692
rect 16206 3680 16212 3732
rect 16264 3720 16270 3732
rect 16301 3723 16359 3729
rect 16301 3720 16313 3723
rect 16264 3692 16313 3720
rect 16264 3680 16270 3692
rect 16301 3689 16313 3692
rect 16347 3689 16359 3723
rect 17494 3720 17500 3732
rect 17455 3692 17500 3720
rect 16301 3683 16359 3689
rect 17494 3680 17500 3692
rect 17552 3680 17558 3732
rect 18141 3723 18199 3729
rect 18141 3689 18153 3723
rect 18187 3720 18199 3723
rect 18414 3720 18420 3732
rect 18187 3692 18420 3720
rect 18187 3689 18199 3692
rect 18141 3683 18199 3689
rect 18414 3680 18420 3692
rect 18472 3680 18478 3732
rect 23106 3720 23112 3732
rect 20180 3692 23112 3720
rect 13998 3612 14004 3664
rect 14056 3652 14062 3664
rect 15473 3655 15531 3661
rect 14056 3624 14964 3652
rect 14056 3612 14062 3624
rect 13354 3544 13360 3596
rect 13412 3584 13418 3596
rect 14826 3584 14832 3596
rect 13412 3556 14832 3584
rect 13412 3544 13418 3556
rect 14826 3544 14832 3556
rect 14884 3544 14890 3596
rect 14936 3584 14964 3624
rect 15473 3621 15485 3655
rect 15519 3652 15531 3655
rect 17034 3652 17040 3664
rect 15519 3624 17040 3652
rect 15519 3621 15531 3624
rect 15473 3615 15531 3621
rect 17034 3612 17040 3624
rect 17092 3612 17098 3664
rect 16945 3587 17003 3593
rect 16945 3584 16957 3587
rect 14936 3556 16957 3584
rect 16945 3553 16957 3556
rect 16991 3584 17003 3587
rect 18785 3587 18843 3593
rect 18785 3584 18797 3587
rect 16991 3556 18797 3584
rect 16991 3553 17003 3556
rect 16945 3547 17003 3553
rect 18785 3553 18797 3556
rect 18831 3584 18843 3587
rect 20180 3584 20208 3692
rect 23106 3680 23112 3692
rect 23164 3680 23170 3732
rect 23382 3680 23388 3732
rect 23440 3720 23446 3732
rect 23753 3723 23811 3729
rect 23753 3720 23765 3723
rect 23440 3692 23765 3720
rect 23440 3680 23446 3692
rect 23753 3689 23765 3692
rect 23799 3689 23811 3723
rect 28074 3720 28080 3732
rect 28035 3692 28080 3720
rect 23753 3683 23811 3689
rect 28074 3680 28080 3692
rect 28132 3680 28138 3732
rect 36722 3720 36728 3732
rect 35866 3692 36728 3720
rect 22465 3655 22523 3661
rect 22465 3621 22477 3655
rect 22511 3621 22523 3655
rect 22465 3615 22523 3621
rect 18831 3556 20208 3584
rect 20257 3587 20315 3593
rect 18831 3553 18843 3556
rect 18785 3547 18843 3553
rect 20257 3553 20269 3587
rect 20303 3584 20315 3587
rect 22002 3584 22008 3596
rect 20303 3556 22008 3584
rect 20303 3553 20315 3556
rect 20257 3547 20315 3553
rect 22002 3544 22008 3556
rect 22060 3544 22066 3596
rect 22186 3544 22192 3596
rect 22244 3584 22250 3596
rect 22480 3584 22508 3615
rect 22554 3612 22560 3664
rect 22612 3652 22618 3664
rect 22612 3624 27108 3652
rect 22612 3612 22618 3624
rect 23106 3584 23112 3596
rect 22244 3556 22508 3584
rect 23067 3556 23112 3584
rect 22244 3544 22250 3556
rect 23106 3544 23112 3556
rect 23164 3544 23170 3596
rect 27080 3584 27108 3624
rect 27154 3612 27160 3664
rect 27212 3652 27218 3664
rect 35866 3652 35894 3692
rect 36722 3680 36728 3692
rect 36780 3680 36786 3732
rect 27212 3624 35894 3652
rect 27212 3612 27218 3624
rect 28902 3584 28908 3596
rect 23952 3556 27016 3584
rect 27080 3556 28396 3584
rect 28863 3556 28908 3584
rect 14550 3476 14556 3528
rect 14608 3516 14614 3528
rect 15013 3519 15071 3525
rect 15013 3516 15025 3519
rect 14608 3488 15025 3516
rect 14608 3476 14614 3488
rect 15013 3485 15025 3488
rect 15059 3485 15071 3519
rect 15013 3479 15071 3485
rect 17681 3519 17739 3525
rect 17681 3485 17693 3519
rect 17727 3516 17739 3519
rect 18046 3516 18052 3528
rect 17727 3488 18052 3516
rect 17727 3485 17739 3488
rect 17681 3479 17739 3485
rect 18046 3476 18052 3488
rect 18104 3476 18110 3528
rect 16761 3451 16819 3457
rect 16761 3448 16773 3451
rect 16546 3420 16773 3448
rect 13219 3352 13308 3380
rect 13219 3349 13231 3352
rect 13173 3343 13231 3349
rect 14550 3340 14556 3392
rect 14608 3380 14614 3392
rect 15105 3383 15163 3389
rect 15105 3380 15117 3383
rect 14608 3352 15117 3380
rect 14608 3340 14614 3352
rect 15105 3349 15117 3352
rect 15151 3380 15163 3383
rect 16546 3380 16574 3420
rect 16761 3417 16773 3420
rect 16807 3417 16819 3451
rect 16761 3411 16819 3417
rect 18509 3451 18567 3457
rect 18509 3417 18521 3451
rect 18555 3448 18567 3451
rect 19794 3448 19800 3460
rect 18555 3420 19800 3448
rect 18555 3417 18567 3420
rect 18509 3411 18567 3417
rect 19794 3408 19800 3420
rect 19852 3408 19858 3460
rect 19886 3408 19892 3460
rect 19944 3448 19950 3460
rect 20533 3451 20591 3457
rect 20533 3448 20545 3451
rect 19944 3420 20545 3448
rect 19944 3408 19950 3420
rect 20533 3417 20545 3420
rect 20579 3417 20591 3451
rect 21910 3448 21916 3460
rect 21758 3420 21916 3448
rect 20533 3411 20591 3417
rect 21910 3408 21916 3420
rect 21968 3408 21974 3460
rect 22020 3448 22048 3544
rect 22833 3519 22891 3525
rect 22833 3485 22845 3519
rect 22879 3516 22891 3519
rect 22922 3516 22928 3528
rect 22879 3488 22928 3516
rect 22879 3485 22891 3488
rect 22833 3479 22891 3485
rect 22922 3476 22928 3488
rect 22980 3476 22986 3528
rect 23842 3516 23848 3528
rect 23755 3488 23848 3516
rect 23842 3476 23848 3488
rect 23900 3516 23906 3528
rect 23952 3516 23980 3556
rect 23900 3488 23980 3516
rect 23900 3476 23906 3488
rect 24578 3476 24584 3528
rect 24636 3516 24642 3528
rect 24765 3519 24823 3525
rect 24765 3516 24777 3519
rect 24636 3488 24777 3516
rect 24636 3476 24642 3488
rect 24765 3485 24777 3488
rect 24811 3516 24823 3519
rect 26988 3516 27016 3556
rect 28368 3528 28396 3556
rect 28902 3544 28908 3556
rect 28960 3544 28966 3596
rect 27985 3519 28043 3525
rect 27985 3516 27997 3519
rect 24811 3488 26234 3516
rect 26988 3488 27997 3516
rect 24811 3485 24823 3488
rect 24765 3479 24823 3485
rect 25038 3448 25044 3460
rect 22020 3420 25044 3448
rect 25038 3408 25044 3420
rect 25096 3408 25102 3460
rect 15151 3352 16574 3380
rect 16669 3383 16727 3389
rect 15151 3349 15163 3352
rect 15105 3343 15163 3349
rect 16669 3349 16681 3383
rect 16715 3380 16727 3383
rect 17862 3380 17868 3392
rect 16715 3352 17868 3380
rect 16715 3349 16727 3352
rect 16669 3343 16727 3349
rect 17862 3340 17868 3352
rect 17920 3340 17926 3392
rect 18598 3340 18604 3392
rect 18656 3380 18662 3392
rect 22002 3380 22008 3392
rect 18656 3352 18701 3380
rect 21963 3352 22008 3380
rect 18656 3340 18662 3352
rect 22002 3340 22008 3352
rect 22060 3380 22066 3392
rect 22925 3383 22983 3389
rect 22925 3380 22937 3383
rect 22060 3352 22937 3380
rect 22060 3340 22066 3352
rect 22925 3349 22937 3352
rect 22971 3349 22983 3383
rect 24670 3380 24676 3392
rect 24631 3352 24676 3380
rect 22925 3343 22983 3349
rect 24670 3340 24676 3352
rect 24728 3340 24734 3392
rect 26206 3380 26234 3488
rect 27985 3485 27997 3488
rect 28031 3485 28043 3519
rect 27985 3479 28043 3485
rect 28000 3448 28028 3479
rect 28350 3476 28356 3528
rect 28408 3516 28414 3528
rect 28629 3519 28687 3525
rect 28629 3516 28641 3519
rect 28408 3488 28641 3516
rect 28408 3476 28414 3488
rect 28629 3485 28641 3488
rect 28675 3485 28687 3519
rect 32766 3516 32772 3528
rect 28629 3479 28687 3485
rect 28828 3488 32772 3516
rect 28828 3448 28856 3488
rect 32766 3476 32772 3488
rect 32824 3476 32830 3528
rect 28000 3420 28856 3448
rect 28902 3380 28908 3392
rect 26206 3352 28908 3380
rect 28902 3340 28908 3352
rect 28960 3340 28966 3392
rect 1104 3290 37628 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 35594 3290
rect 35646 3238 35658 3290
rect 35710 3238 35722 3290
rect 35774 3238 35786 3290
rect 35838 3238 35850 3290
rect 35902 3238 37628 3290
rect 1104 3216 37628 3238
rect 11149 3179 11207 3185
rect 11149 3145 11161 3179
rect 11195 3176 11207 3179
rect 11195 3148 12664 3176
rect 11195 3145 11207 3148
rect 11149 3139 11207 3145
rect 12342 3108 12348 3120
rect 10980 3080 12348 3108
rect 1765 3043 1823 3049
rect 1765 3009 1777 3043
rect 1811 3040 1823 3043
rect 7834 3040 7840 3052
rect 1811 3012 7840 3040
rect 1811 3009 1823 3012
rect 1765 3003 1823 3009
rect 7834 3000 7840 3012
rect 7892 3000 7898 3052
rect 10980 3049 11008 3080
rect 12342 3068 12348 3080
rect 12400 3068 12406 3120
rect 12636 3117 12664 3148
rect 12986 3136 12992 3188
rect 13044 3176 13050 3188
rect 14093 3179 14151 3185
rect 14093 3176 14105 3179
rect 13044 3148 14105 3176
rect 13044 3136 13050 3148
rect 14093 3145 14105 3148
rect 14139 3145 14151 3179
rect 19886 3176 19892 3188
rect 19847 3148 19892 3176
rect 14093 3139 14151 3145
rect 19886 3136 19892 3148
rect 19944 3136 19950 3188
rect 19978 3136 19984 3188
rect 20036 3176 20042 3188
rect 20349 3179 20407 3185
rect 20349 3176 20361 3179
rect 20036 3148 20361 3176
rect 20036 3136 20042 3148
rect 20349 3145 20361 3148
rect 20395 3145 20407 3179
rect 20349 3139 20407 3145
rect 21358 3136 21364 3188
rect 21416 3176 21422 3188
rect 26234 3176 26240 3188
rect 21416 3148 26240 3176
rect 21416 3136 21422 3148
rect 26234 3136 26240 3148
rect 26292 3136 26298 3188
rect 12621 3111 12679 3117
rect 12621 3077 12633 3111
rect 12667 3077 12679 3111
rect 12621 3071 12679 3077
rect 13078 3068 13084 3120
rect 13136 3068 13142 3120
rect 16025 3111 16083 3117
rect 16025 3077 16037 3111
rect 16071 3108 16083 3111
rect 16850 3108 16856 3120
rect 16071 3080 16856 3108
rect 16071 3077 16083 3080
rect 16025 3071 16083 3077
rect 16850 3068 16856 3080
rect 16908 3068 16914 3120
rect 18690 3108 18696 3120
rect 18630 3080 18696 3108
rect 18690 3068 18696 3080
rect 18748 3068 18754 3120
rect 20717 3111 20775 3117
rect 20717 3077 20729 3111
rect 20763 3108 20775 3111
rect 22186 3108 22192 3120
rect 20763 3080 22192 3108
rect 20763 3077 20775 3080
rect 20717 3071 20775 3077
rect 22186 3068 22192 3080
rect 22244 3068 22250 3120
rect 22554 3108 22560 3120
rect 22515 3080 22560 3108
rect 22554 3068 22560 3080
rect 22612 3068 22618 3120
rect 24670 3108 24676 3120
rect 24334 3080 24676 3108
rect 24670 3068 24676 3080
rect 24728 3068 24734 3120
rect 10965 3043 11023 3049
rect 10965 3009 10977 3043
rect 11011 3009 11023 3043
rect 10965 3003 11023 3009
rect 11701 3043 11759 3049
rect 11701 3009 11713 3043
rect 11747 3009 11759 3043
rect 11701 3003 11759 3009
rect 1578 2836 1584 2848
rect 1539 2808 1584 2836
rect 1578 2796 1584 2808
rect 1636 2796 1642 2848
rect 11716 2836 11744 3003
rect 14918 3000 14924 3052
rect 14976 3000 14982 3052
rect 16298 3000 16304 3052
rect 16356 3040 16362 3052
rect 17129 3043 17187 3049
rect 17129 3040 17141 3043
rect 16356 3012 17141 3040
rect 16356 3000 16362 3012
rect 17129 3009 17141 3012
rect 17175 3009 17187 3043
rect 19702 3040 19708 3052
rect 19663 3012 19708 3040
rect 17129 3003 17187 3009
rect 19702 3000 19708 3012
rect 19760 3000 19766 3052
rect 19794 3000 19800 3052
rect 19852 3040 19858 3052
rect 20530 3040 20536 3052
rect 19852 3012 20536 3040
rect 19852 3000 19858 3012
rect 20530 3000 20536 3012
rect 20588 3040 20594 3052
rect 20809 3043 20867 3049
rect 20809 3040 20821 3043
rect 20588 3012 20821 3040
rect 20588 3000 20594 3012
rect 20809 3009 20821 3012
rect 20855 3009 20867 3043
rect 20809 3003 20867 3009
rect 22833 3043 22891 3049
rect 22833 3009 22845 3043
rect 22879 3009 22891 3043
rect 22833 3003 22891 3009
rect 12158 2932 12164 2984
rect 12216 2972 12222 2984
rect 12345 2975 12403 2981
rect 12345 2972 12357 2975
rect 12216 2944 12357 2972
rect 12216 2932 12222 2944
rect 12345 2941 12357 2944
rect 12391 2941 12403 2975
rect 15286 2972 15292 2984
rect 12345 2935 12403 2941
rect 12452 2944 15292 2972
rect 11885 2907 11943 2913
rect 11885 2873 11897 2907
rect 11931 2904 11943 2907
rect 12452 2904 12480 2944
rect 15286 2932 15292 2944
rect 15344 2932 15350 2984
rect 17402 2972 17408 2984
rect 17363 2944 17408 2972
rect 17402 2932 17408 2944
rect 17460 2932 17466 2984
rect 20993 2975 21051 2981
rect 20993 2941 21005 2975
rect 21039 2972 21051 2975
rect 22646 2972 22652 2984
rect 21039 2944 22652 2972
rect 21039 2941 21051 2944
rect 20993 2935 21051 2941
rect 22646 2932 22652 2944
rect 22704 2932 22710 2984
rect 22848 2972 22876 3003
rect 25038 3000 25044 3052
rect 25096 3040 25102 3052
rect 36722 3040 36728 3052
rect 25096 3012 25141 3040
rect 36683 3012 36728 3040
rect 25096 3000 25102 3012
rect 36722 3000 36728 3012
rect 36780 3000 36786 3052
rect 24762 2972 24768 2984
rect 22848 2944 23796 2972
rect 24723 2944 24768 2972
rect 11931 2876 12480 2904
rect 11931 2873 11943 2876
rect 11885 2867 11943 2873
rect 23014 2864 23020 2916
rect 23072 2904 23078 2916
rect 23293 2907 23351 2913
rect 23293 2904 23305 2907
rect 23072 2876 23305 2904
rect 23072 2864 23078 2876
rect 23293 2873 23305 2876
rect 23339 2873 23351 2907
rect 23293 2867 23351 2873
rect 12802 2836 12808 2848
rect 11716 2808 12808 2836
rect 12802 2796 12808 2808
rect 12860 2796 12866 2848
rect 14550 2836 14556 2848
rect 14511 2808 14556 2836
rect 14550 2796 14556 2808
rect 14608 2796 14614 2848
rect 18046 2796 18052 2848
rect 18104 2836 18110 2848
rect 18598 2836 18604 2848
rect 18104 2808 18604 2836
rect 18104 2796 18110 2808
rect 18598 2796 18604 2808
rect 18656 2836 18662 2848
rect 18877 2839 18935 2845
rect 18877 2836 18889 2839
rect 18656 2808 18889 2836
rect 18656 2796 18662 2808
rect 18877 2805 18889 2808
rect 18923 2805 18935 2839
rect 23768 2836 23796 2944
rect 24762 2932 24768 2944
rect 24820 2932 24826 2984
rect 25222 2836 25228 2848
rect 23768 2808 25228 2836
rect 18877 2799 18935 2805
rect 25222 2796 25228 2808
rect 25280 2796 25286 2848
rect 36906 2836 36912 2848
rect 36867 2808 36912 2836
rect 36906 2796 36912 2808
rect 36964 2796 36970 2848
rect 1104 2746 37628 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 37628 2746
rect 1104 2672 37628 2694
rect 10505 2635 10563 2641
rect 10505 2601 10517 2635
rect 10551 2632 10563 2635
rect 12434 2632 12440 2644
rect 10551 2604 12440 2632
rect 10551 2601 10563 2604
rect 10505 2595 10563 2601
rect 12434 2592 12440 2604
rect 12492 2592 12498 2644
rect 14918 2632 14924 2644
rect 14879 2604 14924 2632
rect 14918 2592 14924 2604
rect 14976 2592 14982 2644
rect 15473 2635 15531 2641
rect 15473 2601 15485 2635
rect 15519 2632 15531 2635
rect 16022 2632 16028 2644
rect 15519 2604 16028 2632
rect 15519 2601 15531 2604
rect 15473 2595 15531 2601
rect 16022 2592 16028 2604
rect 16080 2592 16086 2644
rect 16301 2635 16359 2641
rect 16301 2601 16313 2635
rect 16347 2632 16359 2635
rect 17402 2632 17408 2644
rect 16347 2604 17408 2632
rect 16347 2601 16359 2604
rect 16301 2595 16359 2601
rect 17402 2592 17408 2604
rect 17460 2592 17466 2644
rect 18690 2632 18696 2644
rect 18651 2604 18696 2632
rect 18690 2592 18696 2604
rect 18748 2592 18754 2644
rect 19702 2592 19708 2644
rect 19760 2632 19766 2644
rect 20073 2635 20131 2641
rect 20073 2632 20085 2635
rect 19760 2604 20085 2632
rect 19760 2592 19766 2604
rect 20073 2601 20085 2604
rect 20119 2601 20131 2635
rect 20073 2595 20131 2601
rect 21910 2592 21916 2644
rect 21968 2632 21974 2644
rect 22097 2635 22155 2641
rect 22097 2632 22109 2635
rect 21968 2604 22109 2632
rect 21968 2592 21974 2604
rect 22097 2601 22109 2604
rect 22143 2601 22155 2635
rect 24762 2632 24768 2644
rect 24723 2604 24768 2632
rect 22097 2595 22155 2601
rect 24762 2592 24768 2604
rect 24820 2592 24826 2644
rect 25222 2632 25228 2644
rect 25183 2604 25228 2632
rect 25222 2592 25228 2604
rect 25280 2592 25286 2644
rect 27062 2592 27068 2644
rect 27120 2632 27126 2644
rect 32539 2635 32597 2641
rect 32539 2632 32551 2635
rect 27120 2604 32551 2632
rect 27120 2592 27126 2604
rect 32539 2601 32551 2604
rect 32585 2601 32597 2635
rect 32539 2595 32597 2601
rect 34790 2592 34796 2644
rect 34848 2632 34854 2644
rect 34885 2635 34943 2641
rect 34885 2632 34897 2635
rect 34848 2604 34897 2632
rect 34848 2592 34854 2604
rect 34885 2601 34897 2604
rect 34931 2601 34943 2635
rect 34885 2595 34943 2601
rect 10962 2524 10968 2576
rect 11020 2564 11026 2576
rect 11701 2567 11759 2573
rect 11701 2564 11713 2567
rect 11020 2536 11713 2564
rect 11020 2524 11026 2536
rect 11701 2533 11713 2536
rect 11747 2533 11759 2567
rect 11701 2527 11759 2533
rect 17586 2524 17592 2576
rect 17644 2564 17650 2576
rect 24578 2564 24584 2576
rect 17644 2536 19656 2564
rect 17644 2524 17650 2536
rect 1762 2428 1768 2440
rect 1723 2400 1768 2428
rect 1762 2388 1768 2400
rect 1820 2388 1826 2440
rect 4430 2428 4436 2440
rect 4391 2400 4436 2428
rect 4430 2388 4436 2400
rect 4488 2388 4494 2440
rect 7190 2428 7196 2440
rect 7151 2400 7196 2428
rect 7190 2388 7196 2400
rect 7248 2388 7254 2440
rect 9861 2431 9919 2437
rect 9861 2397 9873 2431
rect 9907 2397 9919 2431
rect 9861 2391 9919 2397
rect 10321 2431 10379 2437
rect 10321 2397 10333 2431
rect 10367 2428 10379 2431
rect 10980 2428 11008 2524
rect 12158 2456 12164 2508
rect 12216 2496 12222 2508
rect 13449 2499 13507 2505
rect 13449 2496 13461 2499
rect 12216 2468 13461 2496
rect 12216 2456 12222 2468
rect 13449 2465 13461 2468
rect 13495 2465 13507 2499
rect 13449 2459 13507 2465
rect 13538 2456 13544 2508
rect 13596 2496 13602 2508
rect 17862 2496 17868 2508
rect 13596 2468 17172 2496
rect 17823 2468 17868 2496
rect 13596 2456 13602 2468
rect 11146 2428 11152 2440
rect 10367 2400 11008 2428
rect 11107 2400 11152 2428
rect 10367 2397 10379 2400
rect 10321 2391 10379 2397
rect 1394 2252 1400 2304
rect 1452 2292 1458 2304
rect 1581 2295 1639 2301
rect 1581 2292 1593 2295
rect 1452 2264 1593 2292
rect 1452 2252 1458 2264
rect 1581 2261 1593 2264
rect 1627 2261 1639 2295
rect 1581 2255 1639 2261
rect 4154 2252 4160 2304
rect 4212 2292 4218 2304
rect 4249 2295 4307 2301
rect 4249 2292 4261 2295
rect 4212 2264 4261 2292
rect 4212 2252 4218 2264
rect 4249 2261 4261 2264
rect 4295 2261 4307 2295
rect 4249 2255 4307 2261
rect 6914 2252 6920 2304
rect 6972 2292 6978 2304
rect 7009 2295 7067 2301
rect 7009 2292 7021 2295
rect 6972 2264 7021 2292
rect 6972 2252 6978 2264
rect 7009 2261 7021 2264
rect 7055 2261 7067 2295
rect 9674 2292 9680 2304
rect 9635 2264 9680 2292
rect 7009 2255 7067 2261
rect 9674 2252 9680 2264
rect 9732 2252 9738 2304
rect 9876 2292 9904 2391
rect 11146 2388 11152 2400
rect 11204 2388 11210 2440
rect 14844 2437 14872 2468
rect 14829 2431 14887 2437
rect 14829 2397 14841 2431
rect 14875 2397 14887 2431
rect 14829 2391 14887 2397
rect 15657 2431 15715 2437
rect 15657 2397 15669 2431
rect 15703 2428 15715 2431
rect 15930 2428 15936 2440
rect 15703 2400 15936 2428
rect 15703 2397 15715 2400
rect 15657 2391 15715 2397
rect 15930 2388 15936 2400
rect 15988 2388 15994 2440
rect 16117 2431 16175 2437
rect 16117 2397 16129 2431
rect 16163 2428 16175 2431
rect 17144 2428 17172 2468
rect 17862 2456 17868 2468
rect 17920 2456 17926 2508
rect 18049 2499 18107 2505
rect 18049 2465 18061 2499
rect 18095 2496 18107 2499
rect 18095 2468 19564 2496
rect 18095 2465 18107 2468
rect 18049 2459 18107 2465
rect 17310 2428 17316 2440
rect 16163 2400 16574 2428
rect 17144 2400 17316 2428
rect 16163 2397 16175 2400
rect 16117 2391 16175 2397
rect 11057 2363 11115 2369
rect 11057 2329 11069 2363
rect 11103 2360 11115 2363
rect 11103 2332 12006 2360
rect 11103 2329 11115 2332
rect 11057 2323 11115 2329
rect 12894 2320 12900 2372
rect 12952 2360 12958 2372
rect 13173 2363 13231 2369
rect 13173 2360 13185 2363
rect 12952 2332 13185 2360
rect 12952 2320 12958 2332
rect 13173 2329 13185 2332
rect 13219 2329 13231 2363
rect 13173 2323 13231 2329
rect 11882 2292 11888 2304
rect 9876 2264 11888 2292
rect 11882 2252 11888 2264
rect 11940 2252 11946 2304
rect 16546 2292 16574 2400
rect 17310 2388 17316 2400
rect 17368 2428 17374 2440
rect 18601 2431 18659 2437
rect 18601 2428 18613 2431
rect 17368 2400 18613 2428
rect 17368 2388 17374 2400
rect 18601 2397 18613 2400
rect 18647 2397 18659 2431
rect 18601 2391 18659 2397
rect 17773 2363 17831 2369
rect 17773 2329 17785 2363
rect 17819 2360 17831 2363
rect 18046 2360 18052 2372
rect 17819 2332 18052 2360
rect 17819 2329 17831 2332
rect 17773 2323 17831 2329
rect 18046 2320 18052 2332
rect 18104 2320 18110 2372
rect 19536 2360 19564 2468
rect 19628 2437 19656 2536
rect 22204 2536 24584 2564
rect 20530 2496 20536 2508
rect 20491 2468 20536 2496
rect 20530 2456 20536 2468
rect 20588 2456 20594 2508
rect 20625 2499 20683 2505
rect 20625 2465 20637 2499
rect 20671 2496 20683 2499
rect 22094 2496 22100 2508
rect 20671 2468 22100 2496
rect 20671 2465 20683 2468
rect 20625 2459 20683 2465
rect 19613 2431 19671 2437
rect 19613 2397 19625 2431
rect 19659 2397 19671 2431
rect 20640 2428 20668 2459
rect 22094 2456 22100 2468
rect 22152 2456 22158 2508
rect 21450 2428 21456 2440
rect 19613 2391 19671 2397
rect 19720 2400 20668 2428
rect 21411 2400 21456 2428
rect 19720 2360 19748 2400
rect 21450 2388 21456 2400
rect 21508 2388 21514 2440
rect 22204 2437 22232 2536
rect 24578 2524 24584 2536
rect 24636 2524 24642 2576
rect 22278 2456 22284 2508
rect 22336 2496 22342 2508
rect 22925 2499 22983 2505
rect 22925 2496 22937 2499
rect 22336 2468 22937 2496
rect 22336 2456 22342 2468
rect 22925 2465 22937 2468
rect 22971 2465 22983 2499
rect 22925 2459 22983 2465
rect 23474 2456 23480 2508
rect 23532 2496 23538 2508
rect 23532 2468 25452 2496
rect 23532 2456 23538 2468
rect 22189 2431 22247 2437
rect 22189 2397 22201 2431
rect 22235 2397 22247 2431
rect 22189 2391 22247 2397
rect 23014 2388 23020 2440
rect 23072 2428 23078 2440
rect 25424 2437 25452 2468
rect 30190 2456 30196 2508
rect 30248 2496 30254 2508
rect 30248 2468 35894 2496
rect 30248 2456 30254 2468
rect 23201 2431 23259 2437
rect 23201 2428 23213 2431
rect 23072 2400 23213 2428
rect 23072 2388 23078 2400
rect 23201 2397 23213 2400
rect 23247 2397 23259 2431
rect 24581 2431 24639 2437
rect 24581 2428 24593 2431
rect 23201 2391 23259 2397
rect 23584 2400 24593 2428
rect 22002 2360 22008 2372
rect 19536 2332 19748 2360
rect 20456 2332 22008 2360
rect 20456 2304 20484 2332
rect 22002 2320 22008 2332
rect 22060 2320 22066 2372
rect 22922 2320 22928 2372
rect 22980 2360 22986 2372
rect 23109 2363 23167 2369
rect 23109 2360 23121 2363
rect 22980 2332 23121 2360
rect 22980 2320 22986 2332
rect 23109 2329 23121 2332
rect 23155 2329 23167 2363
rect 23109 2323 23167 2329
rect 17405 2295 17463 2301
rect 17405 2292 17417 2295
rect 16546 2264 17417 2292
rect 17405 2261 17417 2264
rect 17451 2261 17463 2295
rect 17405 2255 17463 2261
rect 17954 2252 17960 2304
rect 18012 2292 18018 2304
rect 19429 2295 19487 2301
rect 19429 2292 19441 2295
rect 18012 2264 19441 2292
rect 18012 2252 18018 2264
rect 19429 2261 19441 2264
rect 19475 2261 19487 2295
rect 20438 2292 20444 2304
rect 20399 2264 20444 2292
rect 19429 2255 19487 2261
rect 20438 2252 20444 2264
rect 20496 2252 20502 2304
rect 20714 2252 20720 2304
rect 20772 2292 20778 2304
rect 23584 2301 23612 2400
rect 24581 2397 24593 2400
rect 24627 2397 24639 2431
rect 24581 2391 24639 2397
rect 25409 2431 25467 2437
rect 25409 2397 25421 2431
rect 25455 2397 25467 2431
rect 25409 2391 25467 2397
rect 31754 2388 31760 2440
rect 31812 2428 31818 2440
rect 32309 2431 32367 2437
rect 32309 2428 32321 2431
rect 31812 2400 32321 2428
rect 31812 2388 31818 2400
rect 32309 2397 32321 2400
rect 32355 2397 32367 2431
rect 32309 2391 32367 2397
rect 34514 2388 34520 2440
rect 34572 2428 34578 2440
rect 35069 2431 35127 2437
rect 35069 2428 35081 2431
rect 34572 2400 35081 2428
rect 34572 2388 34578 2400
rect 35069 2397 35081 2400
rect 35115 2397 35127 2431
rect 35866 2428 35894 2468
rect 36725 2431 36783 2437
rect 36725 2428 36737 2431
rect 35866 2400 36737 2428
rect 35069 2391 35127 2397
rect 36725 2397 36737 2400
rect 36771 2397 36783 2431
rect 36725 2391 36783 2397
rect 24486 2320 24492 2372
rect 24544 2360 24550 2372
rect 24544 2332 26234 2360
rect 24544 2320 24550 2332
rect 21269 2295 21327 2301
rect 21269 2292 21281 2295
rect 20772 2264 21281 2292
rect 20772 2252 20778 2264
rect 21269 2261 21281 2264
rect 21315 2261 21327 2295
rect 21269 2255 21327 2261
rect 23569 2295 23627 2301
rect 23569 2261 23581 2295
rect 23615 2261 23627 2295
rect 26206 2292 26234 2332
rect 28994 2320 29000 2372
rect 29052 2360 29058 2372
rect 29825 2363 29883 2369
rect 29825 2360 29837 2363
rect 29052 2332 29837 2360
rect 29052 2320 29058 2332
rect 29825 2329 29837 2332
rect 29871 2329 29883 2363
rect 29825 2323 29883 2329
rect 29917 2295 29975 2301
rect 29917 2292 29929 2295
rect 26206 2264 29929 2292
rect 23569 2255 23627 2261
rect 29917 2261 29929 2264
rect 29963 2261 29975 2295
rect 29917 2255 29975 2261
rect 36909 2295 36967 2301
rect 36909 2261 36921 2295
rect 36955 2292 36967 2295
rect 37274 2292 37280 2304
rect 36955 2264 37280 2292
rect 36955 2261 36967 2264
rect 36909 2255 36967 2261
rect 37274 2252 37280 2264
rect 37332 2252 37338 2304
rect 1104 2202 37628 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 35594 2202
rect 35646 2150 35658 2202
rect 35710 2150 35722 2202
rect 35774 2150 35786 2202
rect 35838 2150 35850 2202
rect 35902 2150 37628 2202
rect 1104 2128 37628 2150
rect 1762 2048 1768 2100
rect 1820 2088 1826 2100
rect 20438 2088 20444 2100
rect 1820 2060 20444 2088
rect 1820 2048 1826 2060
rect 20438 2048 20444 2060
rect 20496 2048 20502 2100
rect 7190 1980 7196 2032
rect 7248 2020 7254 2032
rect 14550 2020 14556 2032
rect 7248 1992 14556 2020
rect 7248 1980 7254 1992
rect 14550 1980 14556 1992
rect 14608 1980 14614 2032
rect 4430 1912 4436 1964
rect 4488 1952 4494 1964
rect 18046 1952 18052 1964
rect 4488 1924 18052 1952
rect 4488 1912 4494 1924
rect 18046 1912 18052 1924
rect 18104 1912 18110 1964
rect 11146 1844 11152 1896
rect 11204 1884 11210 1896
rect 13538 1884 13544 1896
rect 11204 1856 13544 1884
rect 11204 1844 11210 1856
rect 13538 1844 13544 1856
rect 13596 1844 13602 1896
<< via1 >>
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 1768 38539 1820 38548
rect 1768 38505 1777 38539
rect 1777 38505 1811 38539
rect 1811 38505 1820 38539
rect 1768 38496 1820 38505
rect 4712 38539 4764 38548
rect 4712 38505 4721 38539
rect 4721 38505 4755 38539
rect 4755 38505 4764 38539
rect 4712 38496 4764 38505
rect 7656 38539 7708 38548
rect 7656 38505 7665 38539
rect 7665 38505 7699 38539
rect 7699 38505 7708 38539
rect 7656 38496 7708 38505
rect 10508 38496 10560 38548
rect 13084 38496 13136 38548
rect 16304 38539 16356 38548
rect 16304 38505 16313 38539
rect 16313 38505 16347 38539
rect 16347 38505 16356 38539
rect 16304 38496 16356 38505
rect 22284 38496 22336 38548
rect 25228 38496 25280 38548
rect 19064 38428 19116 38480
rect 30288 38496 30340 38548
rect 34060 38496 34112 38548
rect 36912 38539 36964 38548
rect 36912 38505 36921 38539
rect 36921 38505 36955 38539
rect 36955 38505 36964 38539
rect 36912 38496 36964 38505
rect 18696 38360 18748 38412
rect 19984 38403 20036 38412
rect 19984 38369 19993 38403
rect 19993 38369 20027 38403
rect 20027 38369 20036 38403
rect 19984 38360 20036 38369
rect 20352 38360 20404 38412
rect 4804 38292 4856 38344
rect 8116 38292 8168 38344
rect 10140 38292 10192 38344
rect 10416 38292 10468 38344
rect 13084 38335 13136 38344
rect 13084 38301 13093 38335
rect 13093 38301 13127 38335
rect 13127 38301 13136 38335
rect 13084 38292 13136 38301
rect 14648 38335 14700 38344
rect 12624 38224 12676 38276
rect 14648 38301 14657 38335
rect 14657 38301 14691 38335
rect 14691 38301 14700 38335
rect 14648 38292 14700 38301
rect 15016 38292 15068 38344
rect 15752 38292 15804 38344
rect 15200 38224 15252 38276
rect 12348 38199 12400 38208
rect 12348 38165 12357 38199
rect 12357 38165 12391 38199
rect 12391 38165 12400 38199
rect 12348 38156 12400 38165
rect 14096 38156 14148 38208
rect 17132 38199 17184 38208
rect 17132 38165 17141 38199
rect 17141 38165 17175 38199
rect 17175 38165 17184 38199
rect 17132 38156 17184 38165
rect 19524 38292 19576 38344
rect 22560 38335 22612 38344
rect 18604 38224 18656 38276
rect 22560 38301 22569 38335
rect 22569 38301 22603 38335
rect 22603 38301 22612 38335
rect 22560 38292 22612 38301
rect 23480 38292 23532 38344
rect 28172 38428 28224 38480
rect 29552 38360 29604 38412
rect 23664 38335 23716 38344
rect 23664 38301 23673 38335
rect 23673 38301 23707 38335
rect 23707 38301 23716 38335
rect 24768 38335 24820 38344
rect 23664 38292 23716 38301
rect 24768 38301 24777 38335
rect 24777 38301 24811 38335
rect 24811 38301 24820 38335
rect 24768 38292 24820 38301
rect 25412 38335 25464 38344
rect 25412 38301 25421 38335
rect 25421 38301 25455 38335
rect 25455 38301 25464 38335
rect 25412 38292 25464 38301
rect 28540 38292 28592 38344
rect 23572 38224 23624 38276
rect 29736 38267 29788 38276
rect 29736 38233 29745 38267
rect 29745 38233 29779 38267
rect 29779 38233 29788 38267
rect 29736 38224 29788 38233
rect 31392 38335 31444 38344
rect 31392 38301 31401 38335
rect 31401 38301 31435 38335
rect 31435 38301 31444 38335
rect 31392 38292 31444 38301
rect 33508 38292 33560 38344
rect 34704 38292 34756 38344
rect 18144 38199 18196 38208
rect 18144 38165 18153 38199
rect 18153 38165 18187 38199
rect 18187 38165 18196 38199
rect 18144 38156 18196 38165
rect 19432 38199 19484 38208
rect 19432 38165 19441 38199
rect 19441 38165 19475 38199
rect 19475 38165 19484 38199
rect 19432 38156 19484 38165
rect 19892 38199 19944 38208
rect 19892 38165 19901 38199
rect 19901 38165 19935 38199
rect 19935 38165 19944 38199
rect 19892 38156 19944 38165
rect 21364 38199 21416 38208
rect 21364 38165 21373 38199
rect 21373 38165 21407 38199
rect 21407 38165 21416 38199
rect 21364 38156 21416 38165
rect 23112 38199 23164 38208
rect 23112 38165 23121 38199
rect 23121 38165 23155 38199
rect 23155 38165 23164 38199
rect 23112 38156 23164 38165
rect 23756 38199 23808 38208
rect 23756 38165 23765 38199
rect 23765 38165 23799 38199
rect 23799 38165 23808 38199
rect 23756 38156 23808 38165
rect 24492 38156 24544 38208
rect 25228 38199 25280 38208
rect 25228 38165 25237 38199
rect 25237 38165 25271 38199
rect 25271 38165 25280 38199
rect 25228 38156 25280 38165
rect 27712 38156 27764 38208
rect 28724 38199 28776 38208
rect 28724 38165 28733 38199
rect 28733 38165 28767 38199
rect 28767 38165 28776 38199
rect 28724 38156 28776 38165
rect 29920 38199 29972 38208
rect 29920 38165 29945 38199
rect 29945 38165 29972 38199
rect 30104 38199 30156 38208
rect 29920 38156 29972 38165
rect 30104 38165 30113 38199
rect 30113 38165 30147 38199
rect 30147 38165 30156 38199
rect 30104 38156 30156 38165
rect 31484 38156 31536 38208
rect 32404 38199 32456 38208
rect 32404 38165 32413 38199
rect 32413 38165 32447 38199
rect 32447 38165 32456 38199
rect 32404 38156 32456 38165
rect 33048 38199 33100 38208
rect 33048 38165 33057 38199
rect 33057 38165 33091 38199
rect 33091 38165 33100 38199
rect 33048 38156 33100 38165
rect 4874 38054 4926 38106
rect 4938 38054 4990 38106
rect 5002 38054 5054 38106
rect 5066 38054 5118 38106
rect 5130 38054 5182 38106
rect 35594 38054 35646 38106
rect 35658 38054 35710 38106
rect 35722 38054 35774 38106
rect 35786 38054 35838 38106
rect 35850 38054 35902 38106
rect 1584 37995 1636 38004
rect 1584 37961 1593 37995
rect 1593 37961 1627 37995
rect 1627 37961 1636 37995
rect 1584 37952 1636 37961
rect 4804 37952 4856 38004
rect 8116 37995 8168 38004
rect 8116 37961 8125 37995
rect 8125 37961 8159 37995
rect 8159 37961 8168 37995
rect 8116 37952 8168 37961
rect 10140 37995 10192 38004
rect 10140 37961 10149 37995
rect 10149 37961 10183 37995
rect 10183 37961 10192 37995
rect 10140 37952 10192 37961
rect 13084 37952 13136 38004
rect 15752 37995 15804 38004
rect 15752 37961 15761 37995
rect 15761 37961 15795 37995
rect 15795 37961 15804 37995
rect 15752 37952 15804 37961
rect 18604 37995 18656 38004
rect 18604 37961 18613 37995
rect 18613 37961 18647 37995
rect 18647 37961 18656 37995
rect 18604 37952 18656 37961
rect 19248 37995 19300 38004
rect 19248 37961 19257 37995
rect 19257 37961 19291 37995
rect 19291 37961 19300 37995
rect 19248 37952 19300 37961
rect 17132 37927 17184 37936
rect 1768 37859 1820 37868
rect 1768 37825 1777 37859
rect 1777 37825 1811 37859
rect 1811 37825 1820 37859
rect 1768 37816 1820 37825
rect 8300 37859 8352 37868
rect 8300 37825 8309 37859
rect 8309 37825 8343 37859
rect 8343 37825 8352 37859
rect 8300 37816 8352 37825
rect 9588 37859 9640 37868
rect 9588 37825 9597 37859
rect 9597 37825 9631 37859
rect 9631 37825 9640 37859
rect 9588 37816 9640 37825
rect 10324 37859 10376 37868
rect 10324 37825 10333 37859
rect 10333 37825 10367 37859
rect 10367 37825 10376 37859
rect 10324 37816 10376 37825
rect 10784 37859 10836 37868
rect 10784 37825 10793 37859
rect 10793 37825 10827 37859
rect 10827 37825 10836 37859
rect 10784 37816 10836 37825
rect 11612 37816 11664 37868
rect 12808 37859 12860 37868
rect 12808 37825 12817 37859
rect 12817 37825 12851 37859
rect 12851 37825 12860 37859
rect 12808 37816 12860 37825
rect 13452 37816 13504 37868
rect 14280 37859 14332 37868
rect 14280 37825 14289 37859
rect 14289 37825 14323 37859
rect 14323 37825 14332 37859
rect 14280 37816 14332 37825
rect 17132 37893 17141 37927
rect 17141 37893 17175 37927
rect 17175 37893 17184 37927
rect 17132 37884 17184 37893
rect 19892 37884 19944 37936
rect 22008 37884 22060 37936
rect 23756 37952 23808 38004
rect 22744 37884 22796 37936
rect 24492 37927 24544 37936
rect 24492 37893 24501 37927
rect 24501 37893 24535 37927
rect 24535 37893 24544 37927
rect 24492 37884 24544 37893
rect 29736 37952 29788 38004
rect 15292 37816 15344 37868
rect 18236 37816 18288 37868
rect 19064 37859 19116 37868
rect 19064 37825 19073 37859
rect 19073 37825 19107 37859
rect 19107 37825 19116 37859
rect 19064 37816 19116 37825
rect 21364 37816 21416 37868
rect 24216 37859 24268 37868
rect 14372 37791 14424 37800
rect 14372 37757 14381 37791
rect 14381 37757 14415 37791
rect 14415 37757 14424 37791
rect 14372 37748 14424 37757
rect 14464 37791 14516 37800
rect 14464 37757 14473 37791
rect 14473 37757 14507 37791
rect 14507 37757 14516 37791
rect 16856 37791 16908 37800
rect 14464 37748 14516 37757
rect 16856 37757 16865 37791
rect 16865 37757 16899 37791
rect 16899 37757 16908 37791
rect 16856 37748 16908 37757
rect 20168 37791 20220 37800
rect 20168 37757 20177 37791
rect 20177 37757 20211 37791
rect 20211 37757 20220 37791
rect 20168 37748 20220 37757
rect 20352 37791 20404 37800
rect 20352 37757 20361 37791
rect 20361 37757 20395 37791
rect 20395 37757 20404 37791
rect 20352 37748 20404 37757
rect 24216 37825 24225 37859
rect 24225 37825 24259 37859
rect 24259 37825 24268 37859
rect 24216 37816 24268 37825
rect 26424 37859 26476 37868
rect 26424 37825 26433 37859
rect 26433 37825 26467 37859
rect 26467 37825 26476 37859
rect 26424 37816 26476 37825
rect 27160 37816 27212 37868
rect 28080 37816 28132 37868
rect 23572 37748 23624 37800
rect 14740 37680 14792 37732
rect 29368 37816 29420 37868
rect 29552 37859 29604 37868
rect 29552 37825 29561 37859
rect 29561 37825 29595 37859
rect 29595 37825 29604 37859
rect 29552 37816 29604 37825
rect 9404 37655 9456 37664
rect 9404 37621 9413 37655
rect 9413 37621 9447 37655
rect 9447 37621 9456 37655
rect 9404 37612 9456 37621
rect 10968 37655 11020 37664
rect 10968 37621 10977 37655
rect 10977 37621 11011 37655
rect 11011 37621 11020 37655
rect 10968 37612 11020 37621
rect 19616 37612 19668 37664
rect 25504 37612 25556 37664
rect 26516 37655 26568 37664
rect 26516 37621 26525 37655
rect 26525 37621 26559 37655
rect 26559 37621 26568 37655
rect 26516 37612 26568 37621
rect 27988 37612 28040 37664
rect 28080 37612 28132 37664
rect 28632 37655 28684 37664
rect 28632 37621 28641 37655
rect 28641 37621 28675 37655
rect 28675 37621 28684 37655
rect 28632 37612 28684 37621
rect 29092 37655 29144 37664
rect 29092 37621 29101 37655
rect 29101 37621 29135 37655
rect 29135 37621 29144 37655
rect 29092 37612 29144 37621
rect 33416 37952 33468 38004
rect 34704 37995 34756 38004
rect 34704 37961 34713 37995
rect 34713 37961 34747 37995
rect 34747 37961 34756 37995
rect 34704 37952 34756 37961
rect 31484 37927 31536 37936
rect 31484 37893 31493 37927
rect 31493 37893 31527 37927
rect 31527 37893 31536 37927
rect 31484 37884 31536 37893
rect 33048 37884 33100 37936
rect 34520 37859 34572 37868
rect 34520 37825 34529 37859
rect 34529 37825 34563 37859
rect 34563 37825 34572 37859
rect 34520 37816 34572 37825
rect 31760 37791 31812 37800
rect 31760 37757 31769 37791
rect 31769 37757 31803 37791
rect 31803 37757 31812 37791
rect 33784 37791 33836 37800
rect 31760 37748 31812 37757
rect 30288 37612 30340 37664
rect 33784 37757 33793 37791
rect 33793 37757 33827 37791
rect 33827 37757 33836 37791
rect 33784 37748 33836 37757
rect 34060 37791 34112 37800
rect 34060 37757 34069 37791
rect 34069 37757 34103 37791
rect 34103 37757 34112 37791
rect 34060 37748 34112 37757
rect 34060 37612 34112 37664
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 13452 37451 13504 37460
rect 13452 37417 13461 37451
rect 13461 37417 13495 37451
rect 13495 37417 13504 37451
rect 13452 37408 13504 37417
rect 14648 37408 14700 37460
rect 14740 37408 14792 37460
rect 22560 37408 22612 37460
rect 24768 37408 24820 37460
rect 28080 37408 28132 37460
rect 33784 37408 33836 37460
rect 27712 37383 27764 37392
rect 27712 37349 27721 37383
rect 27721 37349 27755 37383
rect 27755 37349 27764 37383
rect 27712 37340 27764 37349
rect 28816 37340 28868 37392
rect 9404 37315 9456 37324
rect 9404 37281 9413 37315
rect 9413 37281 9447 37315
rect 9447 37281 9456 37315
rect 9404 37272 9456 37281
rect 13820 37272 13872 37324
rect 15108 37315 15160 37324
rect 15108 37281 15117 37315
rect 15117 37281 15151 37315
rect 15151 37281 15160 37315
rect 15108 37272 15160 37281
rect 18696 37272 18748 37324
rect 23572 37272 23624 37324
rect 24216 37272 24268 37324
rect 24860 37272 24912 37324
rect 25228 37315 25280 37324
rect 25228 37281 25237 37315
rect 25237 37281 25271 37315
rect 25271 37281 25280 37315
rect 25228 37272 25280 37281
rect 27988 37272 28040 37324
rect 30012 37315 30064 37324
rect 8116 37204 8168 37256
rect 8208 37136 8260 37188
rect 10876 37111 10928 37120
rect 10876 37077 10885 37111
rect 10885 37077 10919 37111
rect 10919 37077 10928 37111
rect 10876 37068 10928 37077
rect 14372 37204 14424 37256
rect 14924 37247 14976 37256
rect 14924 37213 14933 37247
rect 14933 37213 14967 37247
rect 14967 37213 14976 37247
rect 14924 37204 14976 37213
rect 11980 37179 12032 37188
rect 11980 37145 11989 37179
rect 11989 37145 12023 37179
rect 12023 37145 12032 37179
rect 11980 37136 12032 37145
rect 12256 37068 12308 37120
rect 12348 37068 12400 37120
rect 15384 37068 15436 37120
rect 19432 37204 19484 37256
rect 19616 37247 19668 37256
rect 19616 37213 19625 37247
rect 19625 37213 19659 37247
rect 19659 37213 19668 37247
rect 19616 37204 19668 37213
rect 20260 37247 20312 37256
rect 20260 37213 20269 37247
rect 20269 37213 20303 37247
rect 20303 37213 20312 37247
rect 20260 37204 20312 37213
rect 23020 37204 23072 37256
rect 28632 37204 28684 37256
rect 30012 37281 30021 37315
rect 30021 37281 30055 37315
rect 30055 37281 30064 37315
rect 30012 37272 30064 37281
rect 29276 37204 29328 37256
rect 31300 37272 31352 37324
rect 31760 37272 31812 37324
rect 32404 37204 32456 37256
rect 33416 37247 33468 37256
rect 33416 37213 33425 37247
rect 33425 37213 33459 37247
rect 33459 37213 33468 37247
rect 33416 37204 33468 37213
rect 33508 37247 33560 37256
rect 33508 37213 33517 37247
rect 33517 37213 33551 37247
rect 33551 37213 33560 37247
rect 33508 37204 33560 37213
rect 16028 37179 16080 37188
rect 16028 37145 16037 37179
rect 16037 37145 16071 37179
rect 16071 37145 16080 37179
rect 16028 37136 16080 37145
rect 17040 37136 17092 37188
rect 18328 37136 18380 37188
rect 20168 37136 20220 37188
rect 16856 37068 16908 37120
rect 17316 37068 17368 37120
rect 17960 37068 18012 37120
rect 18604 37068 18656 37120
rect 19708 37068 19760 37120
rect 21272 37136 21324 37188
rect 25504 37136 25556 37188
rect 26516 37136 26568 37188
rect 27988 37179 28040 37188
rect 27988 37145 27997 37179
rect 27997 37145 28031 37179
rect 28031 37145 28040 37179
rect 27988 37136 28040 37145
rect 29092 37136 29144 37188
rect 30380 37136 30432 37188
rect 22008 37111 22060 37120
rect 22008 37077 22017 37111
rect 22017 37077 22051 37111
rect 22051 37077 22060 37111
rect 22008 37068 22060 37077
rect 22376 37068 22428 37120
rect 23664 37111 23716 37120
rect 23664 37077 23673 37111
rect 23673 37077 23707 37111
rect 23707 37077 23716 37111
rect 26700 37111 26752 37120
rect 23664 37068 23716 37077
rect 26700 37077 26709 37111
rect 26709 37077 26743 37111
rect 26743 37077 26752 37111
rect 26700 37068 26752 37077
rect 28816 37111 28868 37120
rect 28816 37077 28825 37111
rect 28825 37077 28859 37111
rect 28859 37077 28868 37111
rect 28816 37068 28868 37077
rect 28908 37111 28960 37120
rect 28908 37077 28917 37111
rect 28917 37077 28951 37111
rect 28951 37077 28960 37111
rect 28908 37068 28960 37077
rect 29368 37068 29420 37120
rect 29828 37068 29880 37120
rect 4874 36966 4926 37018
rect 4938 36966 4990 37018
rect 5002 36966 5054 37018
rect 5066 36966 5118 37018
rect 5130 36966 5182 37018
rect 35594 36966 35646 37018
rect 35658 36966 35710 37018
rect 35722 36966 35774 37018
rect 35786 36966 35838 37018
rect 35850 36966 35902 37018
rect 8300 36864 8352 36916
rect 11980 36864 12032 36916
rect 10232 36796 10284 36848
rect 13452 36864 13504 36916
rect 14924 36864 14976 36916
rect 16028 36864 16080 36916
rect 9404 36728 9456 36780
rect 9956 36660 10008 36712
rect 10876 36728 10928 36780
rect 11244 36728 11296 36780
rect 10600 36660 10652 36712
rect 8116 36592 8168 36644
rect 12624 36660 12676 36712
rect 13084 36703 13136 36712
rect 13084 36669 13093 36703
rect 13093 36669 13127 36703
rect 13127 36669 13136 36703
rect 13084 36660 13136 36669
rect 13820 36796 13872 36848
rect 14096 36839 14148 36848
rect 14096 36805 14105 36839
rect 14105 36805 14139 36839
rect 14139 36805 14148 36839
rect 14096 36796 14148 36805
rect 15200 36728 15252 36780
rect 17960 36864 18012 36916
rect 18328 36864 18380 36916
rect 19156 36796 19208 36848
rect 21272 36864 21324 36916
rect 23664 36864 23716 36916
rect 24400 36864 24452 36916
rect 31392 36864 31444 36916
rect 19708 36796 19760 36848
rect 22376 36839 22428 36848
rect 18328 36728 18380 36780
rect 22376 36805 22385 36839
rect 22385 36805 22419 36839
rect 22419 36805 22428 36839
rect 22376 36796 22428 36805
rect 23112 36796 23164 36848
rect 26700 36796 26752 36848
rect 27988 36839 28040 36848
rect 21272 36771 21324 36780
rect 21272 36737 21281 36771
rect 21281 36737 21315 36771
rect 21315 36737 21324 36771
rect 21272 36728 21324 36737
rect 13820 36703 13872 36712
rect 13820 36669 13829 36703
rect 13829 36669 13863 36703
rect 13863 36669 13872 36703
rect 13820 36660 13872 36669
rect 15108 36660 15160 36712
rect 17132 36660 17184 36712
rect 9128 36567 9180 36576
rect 9128 36533 9137 36567
rect 9137 36533 9171 36567
rect 9171 36533 9180 36567
rect 9128 36524 9180 36533
rect 12072 36524 12124 36576
rect 19432 36524 19484 36576
rect 20260 36660 20312 36712
rect 22100 36703 22152 36712
rect 22100 36669 22109 36703
rect 22109 36669 22143 36703
rect 22143 36669 22152 36703
rect 22100 36660 22152 36669
rect 23480 36524 23532 36576
rect 25504 36728 25556 36780
rect 26148 36728 26200 36780
rect 27988 36805 27997 36839
rect 27997 36805 28031 36839
rect 28031 36805 28040 36839
rect 27988 36796 28040 36805
rect 28540 36796 28592 36848
rect 34060 36839 34112 36848
rect 24032 36524 24084 36576
rect 24952 36660 25004 36712
rect 25412 36592 25464 36644
rect 34060 36805 34069 36839
rect 34069 36805 34103 36839
rect 34103 36805 34112 36839
rect 34060 36796 34112 36805
rect 29828 36771 29880 36780
rect 29828 36737 29837 36771
rect 29837 36737 29871 36771
rect 29871 36737 29880 36771
rect 29828 36728 29880 36737
rect 30288 36728 30340 36780
rect 33600 36728 33652 36780
rect 30104 36660 30156 36712
rect 30380 36660 30432 36712
rect 30012 36592 30064 36644
rect 27252 36567 27304 36576
rect 27252 36533 27261 36567
rect 27261 36533 27295 36567
rect 27295 36533 27304 36567
rect 27252 36524 27304 36533
rect 28172 36524 28224 36576
rect 29092 36524 29144 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 9588 36363 9640 36372
rect 9588 36329 9597 36363
rect 9597 36329 9631 36363
rect 9631 36329 9640 36363
rect 9588 36320 9640 36329
rect 9404 36252 9456 36304
rect 11244 36320 11296 36372
rect 17040 36320 17092 36372
rect 18144 36363 18196 36372
rect 18144 36329 18153 36363
rect 18153 36329 18187 36363
rect 18187 36329 18196 36363
rect 18144 36320 18196 36329
rect 22744 36320 22796 36372
rect 23020 36363 23072 36372
rect 23020 36329 23029 36363
rect 23029 36329 23063 36363
rect 23063 36329 23072 36363
rect 23020 36320 23072 36329
rect 12256 36252 12308 36304
rect 13820 36252 13872 36304
rect 18236 36252 18288 36304
rect 18604 36252 18656 36304
rect 27160 36320 27212 36372
rect 30288 36320 30340 36372
rect 31208 36320 31260 36372
rect 8024 36184 8076 36236
rect 12440 36184 12492 36236
rect 13452 36227 13504 36236
rect 13452 36193 13461 36227
rect 13461 36193 13495 36227
rect 13495 36193 13504 36227
rect 13452 36184 13504 36193
rect 16028 36184 16080 36236
rect 19708 36184 19760 36236
rect 19984 36184 20036 36236
rect 23480 36227 23532 36236
rect 23480 36193 23489 36227
rect 23489 36193 23523 36227
rect 23523 36193 23532 36227
rect 23480 36184 23532 36193
rect 23572 36227 23624 36236
rect 23572 36193 23581 36227
rect 23581 36193 23615 36227
rect 23615 36193 23624 36227
rect 23572 36184 23624 36193
rect 24952 36184 25004 36236
rect 7104 36116 7156 36168
rect 8116 36116 8168 36168
rect 9956 36159 10008 36168
rect 9956 36125 9965 36159
rect 9965 36125 9999 36159
rect 9999 36125 10008 36159
rect 9956 36116 10008 36125
rect 10416 36116 10468 36168
rect 13084 36116 13136 36168
rect 17040 36159 17092 36168
rect 17040 36125 17049 36159
rect 17049 36125 17083 36159
rect 17083 36125 17092 36159
rect 17040 36116 17092 36125
rect 17684 36159 17736 36168
rect 17684 36125 17693 36159
rect 17693 36125 17727 36159
rect 17727 36125 17736 36159
rect 17684 36116 17736 36125
rect 17960 36116 18012 36168
rect 18328 36116 18380 36168
rect 19524 36116 19576 36168
rect 20168 36116 20220 36168
rect 27620 36184 27672 36236
rect 29000 36252 29052 36304
rect 31300 36227 31352 36236
rect 31300 36193 31309 36227
rect 31309 36193 31343 36227
rect 31343 36193 31352 36227
rect 31300 36184 31352 36193
rect 32312 36184 32364 36236
rect 26424 36159 26476 36168
rect 10968 36048 11020 36100
rect 12072 36048 12124 36100
rect 7380 35980 7432 36032
rect 7472 35980 7524 36032
rect 8116 35980 8168 36032
rect 8300 36023 8352 36032
rect 8300 35989 8309 36023
rect 8309 35989 8343 36023
rect 8343 35989 8352 36023
rect 8300 35980 8352 35989
rect 10692 35980 10744 36032
rect 14924 36048 14976 36100
rect 17316 36048 17368 36100
rect 19432 36048 19484 36100
rect 21272 36048 21324 36100
rect 26424 36125 26433 36159
rect 26433 36125 26467 36159
rect 26467 36125 26476 36159
rect 26424 36116 26476 36125
rect 27988 36116 28040 36168
rect 30564 36116 30616 36168
rect 30840 36159 30892 36168
rect 30840 36125 30849 36159
rect 30849 36125 30883 36159
rect 30883 36125 30892 36159
rect 30840 36116 30892 36125
rect 33508 36116 33560 36168
rect 26976 36048 27028 36100
rect 28448 36048 28500 36100
rect 30288 36048 30340 36100
rect 33048 36048 33100 36100
rect 12992 36023 13044 36032
rect 12992 35989 13001 36023
rect 13001 35989 13035 36023
rect 13035 35989 13044 36023
rect 12992 35980 13044 35989
rect 15568 36023 15620 36032
rect 15568 35989 15577 36023
rect 15577 35989 15611 36023
rect 15611 35989 15620 36023
rect 15568 35980 15620 35989
rect 19984 36023 20036 36032
rect 19984 35989 19993 36023
rect 19993 35989 20027 36023
rect 20027 35989 20036 36023
rect 19984 35980 20036 35989
rect 20444 36023 20496 36032
rect 20444 35989 20453 36023
rect 20453 35989 20487 36023
rect 20487 35989 20496 36023
rect 20444 35980 20496 35989
rect 23388 36023 23440 36032
rect 23388 35989 23397 36023
rect 23397 35989 23431 36023
rect 23431 35989 23440 36023
rect 23388 35980 23440 35989
rect 24952 36023 25004 36032
rect 24952 35989 24961 36023
rect 24961 35989 24995 36023
rect 24995 35989 25004 36023
rect 24952 35980 25004 35989
rect 25136 35980 25188 36032
rect 26516 36023 26568 36032
rect 26516 35989 26525 36023
rect 26525 35989 26559 36023
rect 26559 35989 26568 36023
rect 26516 35980 26568 35989
rect 28264 35980 28316 36032
rect 28540 36023 28592 36032
rect 28540 35989 28549 36023
rect 28549 35989 28583 36023
rect 28583 35989 28592 36023
rect 28540 35980 28592 35989
rect 29736 36023 29788 36032
rect 29736 35989 29745 36023
rect 29745 35989 29779 36023
rect 29779 35989 29788 36023
rect 29736 35980 29788 35989
rect 31668 35980 31720 36032
rect 33692 35980 33744 36032
rect 4874 35878 4926 35930
rect 4938 35878 4990 35930
rect 5002 35878 5054 35930
rect 5066 35878 5118 35930
rect 5130 35878 5182 35930
rect 35594 35878 35646 35930
rect 35658 35878 35710 35930
rect 35722 35878 35774 35930
rect 35786 35878 35838 35930
rect 35850 35878 35902 35930
rect 10692 35819 10744 35828
rect 10692 35785 10701 35819
rect 10701 35785 10735 35819
rect 10735 35785 10744 35819
rect 10692 35776 10744 35785
rect 10784 35776 10836 35828
rect 12992 35776 13044 35828
rect 7472 35708 7524 35760
rect 7196 35683 7248 35692
rect 7196 35649 7205 35683
rect 7205 35649 7239 35683
rect 7239 35649 7248 35683
rect 7196 35640 7248 35649
rect 8208 35708 8260 35760
rect 9128 35708 9180 35760
rect 9956 35708 10008 35760
rect 15568 35776 15620 35828
rect 19156 35819 19208 35828
rect 19156 35785 19165 35819
rect 19165 35785 19199 35819
rect 19199 35785 19208 35819
rect 19156 35776 19208 35785
rect 20444 35776 20496 35828
rect 23388 35776 23440 35828
rect 24952 35776 25004 35828
rect 14280 35683 14332 35692
rect 10692 35572 10744 35624
rect 6736 35479 6788 35488
rect 6736 35445 6745 35479
rect 6745 35445 6779 35479
rect 6779 35445 6788 35479
rect 6736 35436 6788 35445
rect 8300 35436 8352 35488
rect 9588 35479 9640 35488
rect 9588 35445 9597 35479
rect 9597 35445 9631 35479
rect 9631 35445 9640 35479
rect 14280 35649 14289 35683
rect 14289 35649 14323 35683
rect 14323 35649 14332 35683
rect 14280 35640 14332 35649
rect 15384 35683 15436 35692
rect 15384 35649 15393 35683
rect 15393 35649 15427 35683
rect 15427 35649 15436 35683
rect 15384 35640 15436 35649
rect 15936 35640 15988 35692
rect 17684 35708 17736 35760
rect 19892 35708 19944 35760
rect 22376 35708 22428 35760
rect 25136 35751 25188 35760
rect 25136 35717 25145 35751
rect 25145 35717 25179 35751
rect 25179 35717 25188 35751
rect 25136 35708 25188 35717
rect 26516 35708 26568 35760
rect 28448 35708 28500 35760
rect 28816 35751 28868 35760
rect 28816 35717 28825 35751
rect 28825 35717 28859 35751
rect 28859 35717 28868 35751
rect 28816 35708 28868 35717
rect 29000 35708 29052 35760
rect 29920 35708 29972 35760
rect 30380 35708 30432 35760
rect 17868 35683 17920 35692
rect 17868 35649 17877 35683
rect 17877 35649 17911 35683
rect 17911 35649 17920 35683
rect 17868 35640 17920 35649
rect 19248 35683 19300 35692
rect 19248 35649 19257 35683
rect 19257 35649 19291 35683
rect 19291 35649 19300 35683
rect 19248 35640 19300 35649
rect 12164 35572 12216 35624
rect 13176 35615 13228 35624
rect 13176 35581 13185 35615
rect 13185 35581 13219 35615
rect 13219 35581 13228 35615
rect 13176 35572 13228 35581
rect 13912 35572 13964 35624
rect 15108 35572 15160 35624
rect 17960 35615 18012 35624
rect 17960 35581 17969 35615
rect 17969 35581 18003 35615
rect 18003 35581 18012 35615
rect 17960 35572 18012 35581
rect 18696 35572 18748 35624
rect 19524 35572 19576 35624
rect 13544 35504 13596 35556
rect 21364 35640 21416 35692
rect 23296 35640 23348 35692
rect 24860 35683 24912 35692
rect 24860 35649 24869 35683
rect 24869 35649 24903 35683
rect 24903 35649 24912 35683
rect 24860 35640 24912 35649
rect 28080 35683 28132 35692
rect 28080 35649 28089 35683
rect 28089 35649 28123 35683
rect 28123 35649 28132 35683
rect 28080 35640 28132 35649
rect 28908 35640 28960 35692
rect 23756 35572 23808 35624
rect 24032 35615 24084 35624
rect 24032 35581 24041 35615
rect 24041 35581 24075 35615
rect 24075 35581 24084 35615
rect 24032 35572 24084 35581
rect 27712 35615 27764 35624
rect 27712 35581 27721 35615
rect 27721 35581 27755 35615
rect 27755 35581 27764 35615
rect 27712 35572 27764 35581
rect 29000 35572 29052 35624
rect 29736 35572 29788 35624
rect 31208 35708 31260 35760
rect 30840 35683 30892 35692
rect 30840 35649 30849 35683
rect 30849 35649 30883 35683
rect 30883 35649 30892 35683
rect 30840 35640 30892 35649
rect 32312 35683 32364 35692
rect 28632 35504 28684 35556
rect 30564 35572 30616 35624
rect 14464 35479 14516 35488
rect 9588 35436 9640 35445
rect 14464 35445 14473 35479
rect 14473 35445 14507 35479
rect 14507 35445 14516 35479
rect 14464 35436 14516 35445
rect 16120 35479 16172 35488
rect 16120 35445 16129 35479
rect 16129 35445 16163 35479
rect 16163 35445 16172 35479
rect 16120 35436 16172 35445
rect 16396 35436 16448 35488
rect 20904 35436 20956 35488
rect 22008 35436 22060 35488
rect 22744 35479 22796 35488
rect 22744 35445 22753 35479
rect 22753 35445 22787 35479
rect 22787 35445 22796 35479
rect 22744 35436 22796 35445
rect 28356 35479 28408 35488
rect 28356 35445 28365 35479
rect 28365 35445 28399 35479
rect 28399 35445 28408 35479
rect 28356 35436 28408 35445
rect 29368 35436 29420 35488
rect 30932 35572 30984 35624
rect 32312 35649 32321 35683
rect 32321 35649 32355 35683
rect 32355 35649 32364 35683
rect 32312 35640 32364 35649
rect 33692 35640 33744 35692
rect 30104 35436 30156 35488
rect 31484 35436 31536 35488
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 6736 35232 6788 35284
rect 8116 35232 8168 35284
rect 10324 35275 10376 35284
rect 8208 35096 8260 35148
rect 10324 35241 10333 35275
rect 10333 35241 10367 35275
rect 10367 35241 10376 35275
rect 10324 35232 10376 35241
rect 17960 35232 18012 35284
rect 12164 35164 12216 35216
rect 2044 35028 2096 35080
rect 10324 35096 10376 35148
rect 10600 35096 10652 35148
rect 10968 35139 11020 35148
rect 10968 35105 10977 35139
rect 10977 35105 11011 35139
rect 11011 35105 11020 35139
rect 10968 35096 11020 35105
rect 13820 35096 13872 35148
rect 14556 35096 14608 35148
rect 16764 35096 16816 35148
rect 17316 35096 17368 35148
rect 19892 35139 19944 35148
rect 19892 35105 19901 35139
rect 19901 35105 19935 35139
rect 19935 35105 19944 35139
rect 19892 35096 19944 35105
rect 19984 35139 20036 35148
rect 19984 35105 19993 35139
rect 19993 35105 20027 35139
rect 20027 35105 20036 35139
rect 19984 35096 20036 35105
rect 20352 35096 20404 35148
rect 12164 35028 12216 35080
rect 7380 34960 7432 35012
rect 11244 34960 11296 35012
rect 12440 35028 12492 35080
rect 12624 35028 12676 35080
rect 13544 35071 13596 35080
rect 13544 35037 13553 35071
rect 13553 35037 13587 35071
rect 13587 35037 13596 35071
rect 13544 35028 13596 35037
rect 19248 35028 19300 35080
rect 21364 35232 21416 35284
rect 22376 35275 22428 35284
rect 22376 35241 22385 35275
rect 22385 35241 22419 35275
rect 22419 35241 22428 35275
rect 22376 35232 22428 35241
rect 23296 35275 23348 35284
rect 23296 35241 23305 35275
rect 23305 35241 23339 35275
rect 23339 35241 23348 35275
rect 23296 35232 23348 35241
rect 27620 35232 27672 35284
rect 28172 35275 28224 35284
rect 28172 35241 28181 35275
rect 28181 35241 28215 35275
rect 28215 35241 28224 35275
rect 28172 35232 28224 35241
rect 28540 35232 28592 35284
rect 28816 35232 28868 35284
rect 29920 35275 29972 35284
rect 29920 35241 29929 35275
rect 29929 35241 29963 35275
rect 29963 35241 29972 35275
rect 29920 35232 29972 35241
rect 33048 35232 33100 35284
rect 22192 35164 22244 35216
rect 26976 35164 27028 35216
rect 22100 35096 22152 35148
rect 23388 35096 23440 35148
rect 23572 35096 23624 35148
rect 25044 35096 25096 35148
rect 26056 35096 26108 35148
rect 22008 35028 22060 35080
rect 26700 35028 26752 35080
rect 27252 35096 27304 35148
rect 28264 35139 28316 35148
rect 27896 35071 27948 35080
rect 27896 35037 27905 35071
rect 27905 35037 27939 35071
rect 27939 35037 27948 35071
rect 27896 35028 27948 35037
rect 28264 35105 28273 35139
rect 28273 35105 28307 35139
rect 28307 35105 28316 35139
rect 28264 35096 28316 35105
rect 32312 35096 32364 35148
rect 13452 34960 13504 35012
rect 1584 34935 1636 34944
rect 1584 34901 1593 34935
rect 1593 34901 1627 34935
rect 1627 34901 1636 34935
rect 1584 34892 1636 34901
rect 8852 34892 8904 34944
rect 9496 34935 9548 34944
rect 9496 34901 9505 34935
rect 9505 34901 9539 34935
rect 9539 34901 9548 34935
rect 9496 34892 9548 34901
rect 10600 34892 10652 34944
rect 11796 34935 11848 34944
rect 11796 34901 11805 34935
rect 11805 34901 11839 34935
rect 11839 34901 11848 34935
rect 11796 34892 11848 34901
rect 12348 34935 12400 34944
rect 12348 34901 12357 34935
rect 12357 34901 12391 34935
rect 12391 34901 12400 34935
rect 12348 34892 12400 34901
rect 12992 34935 13044 34944
rect 12992 34901 13001 34935
rect 13001 34901 13035 34935
rect 13035 34901 13044 34935
rect 12992 34892 13044 34901
rect 15568 34960 15620 35012
rect 16304 34960 16356 35012
rect 19524 34960 19576 35012
rect 20904 35003 20956 35012
rect 15936 34892 15988 34944
rect 19340 34892 19392 34944
rect 19800 34935 19852 34944
rect 19800 34901 19809 34935
rect 19809 34901 19843 34935
rect 19843 34901 19852 34935
rect 19800 34892 19852 34901
rect 20904 34969 20913 35003
rect 20913 34969 20947 35003
rect 20947 34969 20956 35003
rect 20904 34960 20956 34969
rect 26148 35003 26200 35012
rect 23388 34892 23440 34944
rect 23940 34892 23992 34944
rect 25688 34892 25740 34944
rect 26148 34969 26157 35003
rect 26157 34969 26191 35003
rect 26191 34969 26200 35003
rect 26148 34960 26200 34969
rect 28448 35028 28500 35080
rect 33508 35028 33560 35080
rect 36912 35071 36964 35080
rect 36912 35037 36921 35071
rect 36921 35037 36955 35071
rect 36955 35037 36964 35071
rect 36912 35028 36964 35037
rect 28540 34960 28592 35012
rect 32680 35003 32732 35012
rect 28264 34892 28316 34944
rect 28448 34892 28500 34944
rect 30564 34892 30616 34944
rect 32680 34969 32689 35003
rect 32689 34969 32723 35003
rect 32723 34969 32732 35003
rect 32680 34960 32732 34969
rect 33140 34892 33192 34944
rect 37096 34935 37148 34944
rect 37096 34901 37105 34935
rect 37105 34901 37139 34935
rect 37139 34901 37148 34935
rect 37096 34892 37148 34901
rect 4874 34790 4926 34842
rect 4938 34790 4990 34842
rect 5002 34790 5054 34842
rect 5066 34790 5118 34842
rect 5130 34790 5182 34842
rect 35594 34790 35646 34842
rect 35658 34790 35710 34842
rect 35722 34790 35774 34842
rect 35786 34790 35838 34842
rect 35850 34790 35902 34842
rect 7196 34688 7248 34740
rect 8852 34731 8904 34740
rect 8852 34697 8861 34731
rect 8861 34697 8895 34731
rect 8895 34697 8904 34731
rect 8852 34688 8904 34697
rect 9588 34688 9640 34740
rect 13176 34688 13228 34740
rect 13452 34688 13504 34740
rect 15568 34731 15620 34740
rect 12348 34620 12400 34672
rect 14556 34620 14608 34672
rect 15568 34697 15577 34731
rect 15577 34697 15611 34731
rect 15611 34697 15620 34731
rect 15568 34688 15620 34697
rect 16304 34731 16356 34740
rect 16304 34697 16313 34731
rect 16313 34697 16347 34731
rect 16347 34697 16356 34731
rect 16304 34688 16356 34697
rect 17868 34688 17920 34740
rect 18604 34688 18656 34740
rect 23940 34731 23992 34740
rect 23940 34697 23949 34731
rect 23949 34697 23983 34731
rect 23983 34697 23992 34731
rect 23940 34688 23992 34697
rect 24952 34688 25004 34740
rect 28264 34731 28316 34740
rect 11244 34552 11296 34604
rect 12072 34595 12124 34604
rect 12072 34561 12081 34595
rect 12081 34561 12115 34595
rect 12115 34561 12124 34595
rect 12072 34552 12124 34561
rect 16396 34552 16448 34604
rect 22744 34620 22796 34672
rect 28264 34697 28273 34731
rect 28273 34697 28307 34731
rect 28307 34697 28316 34731
rect 28264 34688 28316 34697
rect 28632 34731 28684 34740
rect 28632 34697 28641 34731
rect 28641 34697 28675 34731
rect 28675 34697 28684 34731
rect 28632 34688 28684 34697
rect 29920 34688 29972 34740
rect 30932 34731 30984 34740
rect 30932 34697 30934 34731
rect 30934 34697 30968 34731
rect 30968 34697 30984 34731
rect 30932 34688 30984 34697
rect 32680 34688 32732 34740
rect 28448 34620 28500 34672
rect 18052 34552 18104 34604
rect 18420 34595 18472 34604
rect 18420 34561 18429 34595
rect 18429 34561 18463 34595
rect 18463 34561 18472 34595
rect 18420 34552 18472 34561
rect 19432 34595 19484 34604
rect 19432 34561 19441 34595
rect 19441 34561 19475 34595
rect 19475 34561 19484 34595
rect 19432 34552 19484 34561
rect 20812 34552 20864 34604
rect 23756 34552 23808 34604
rect 25688 34552 25740 34604
rect 27252 34552 27304 34604
rect 29000 34552 29052 34604
rect 31116 34620 31168 34672
rect 29920 34595 29972 34604
rect 29920 34561 29929 34595
rect 29929 34561 29963 34595
rect 29963 34561 29972 34595
rect 29920 34552 29972 34561
rect 10692 34484 10744 34536
rect 11152 34484 11204 34536
rect 11980 34484 12032 34536
rect 9680 34416 9732 34468
rect 10876 34416 10928 34468
rect 13912 34484 13964 34536
rect 16028 34416 16080 34468
rect 19800 34484 19852 34536
rect 22100 34484 22152 34536
rect 23940 34484 23992 34536
rect 26056 34484 26108 34536
rect 29460 34484 29512 34536
rect 30380 34484 30432 34536
rect 30472 34484 30524 34536
rect 31208 34552 31260 34604
rect 31484 34595 31536 34604
rect 31484 34561 31493 34595
rect 31493 34561 31527 34595
rect 31527 34561 31536 34595
rect 31484 34552 31536 34561
rect 31668 34595 31720 34604
rect 31668 34561 31677 34595
rect 31677 34561 31711 34595
rect 31711 34561 31720 34595
rect 31668 34552 31720 34561
rect 10692 34348 10744 34400
rect 16120 34348 16172 34400
rect 17868 34348 17920 34400
rect 18236 34348 18288 34400
rect 24860 34416 24912 34468
rect 30288 34459 30340 34468
rect 30288 34425 30297 34459
rect 30297 34425 30331 34459
rect 30331 34425 30340 34459
rect 30288 34416 30340 34425
rect 33600 34459 33652 34468
rect 33600 34425 33609 34459
rect 33609 34425 33643 34459
rect 33643 34425 33652 34459
rect 33600 34416 33652 34425
rect 22192 34348 22244 34400
rect 24400 34391 24452 34400
rect 24400 34357 24409 34391
rect 24409 34357 24443 34391
rect 24443 34357 24452 34391
rect 24400 34348 24452 34357
rect 26240 34391 26292 34400
rect 26240 34357 26249 34391
rect 26249 34357 26283 34391
rect 26283 34357 26292 34391
rect 26240 34348 26292 34357
rect 27896 34348 27948 34400
rect 28632 34348 28684 34400
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 12164 34144 12216 34196
rect 15292 34144 15344 34196
rect 18236 34187 18288 34196
rect 18236 34153 18245 34187
rect 18245 34153 18279 34187
rect 18279 34153 18288 34187
rect 18236 34144 18288 34153
rect 20812 34187 20864 34196
rect 17040 34076 17092 34128
rect 20812 34153 20821 34187
rect 20821 34153 20855 34187
rect 20855 34153 20864 34187
rect 20812 34144 20864 34153
rect 26700 34187 26752 34196
rect 26700 34153 26709 34187
rect 26709 34153 26743 34187
rect 26743 34153 26752 34187
rect 26700 34144 26752 34153
rect 27712 34144 27764 34196
rect 33140 34187 33192 34196
rect 33140 34153 33149 34187
rect 33149 34153 33183 34187
rect 33183 34153 33192 34187
rect 33140 34144 33192 34153
rect 8024 34008 8076 34060
rect 9496 34008 9548 34060
rect 9680 34051 9732 34060
rect 9680 34017 9689 34051
rect 9689 34017 9723 34051
rect 9723 34017 9732 34051
rect 10692 34051 10744 34060
rect 9680 34008 9732 34017
rect 10692 34017 10701 34051
rect 10701 34017 10735 34051
rect 10735 34017 10744 34051
rect 10692 34008 10744 34017
rect 12532 34008 12584 34060
rect 14188 34008 14240 34060
rect 14648 34008 14700 34060
rect 16028 34008 16080 34060
rect 8208 33940 8260 33992
rect 9772 33940 9824 33992
rect 10416 33983 10468 33992
rect 10416 33949 10425 33983
rect 10425 33949 10459 33983
rect 10459 33949 10468 33983
rect 10416 33940 10468 33949
rect 7380 33804 7432 33856
rect 8484 33872 8536 33924
rect 9588 33872 9640 33924
rect 11152 33872 11204 33924
rect 15936 33983 15988 33992
rect 15936 33949 15945 33983
rect 15945 33949 15979 33983
rect 15979 33949 15988 33983
rect 15936 33940 15988 33949
rect 17408 33983 17460 33992
rect 17408 33949 17417 33983
rect 17417 33949 17451 33983
rect 17451 33949 17460 33983
rect 17408 33940 17460 33949
rect 19340 34008 19392 34060
rect 19984 34008 20036 34060
rect 23388 34051 23440 34060
rect 23388 34017 23397 34051
rect 23397 34017 23431 34051
rect 23431 34017 23440 34051
rect 23388 34008 23440 34017
rect 24860 34008 24912 34060
rect 26240 34008 26292 34060
rect 20904 33983 20956 33992
rect 20904 33949 20913 33983
rect 20913 33949 20947 33983
rect 20947 33949 20956 33983
rect 20904 33940 20956 33949
rect 21272 33940 21324 33992
rect 21364 33940 21416 33992
rect 24400 33940 24452 33992
rect 28264 34076 28316 34128
rect 9128 33847 9180 33856
rect 9128 33813 9137 33847
rect 9137 33813 9171 33847
rect 9171 33813 9180 33847
rect 9128 33804 9180 33813
rect 9496 33847 9548 33856
rect 9496 33813 9505 33847
rect 9505 33813 9539 33847
rect 9539 33813 9548 33847
rect 9496 33804 9548 33813
rect 11980 33804 12032 33856
rect 12164 33847 12216 33856
rect 12164 33813 12173 33847
rect 12173 33813 12207 33847
rect 12207 33813 12216 33847
rect 12164 33804 12216 33813
rect 12900 33804 12952 33856
rect 19064 33872 19116 33924
rect 26608 33872 26660 33924
rect 28172 33940 28224 33992
rect 28540 33940 28592 33992
rect 28632 33940 28684 33992
rect 30472 33940 30524 33992
rect 32772 33940 32824 33992
rect 33508 33940 33560 33992
rect 28448 33872 28500 33924
rect 13912 33804 13964 33856
rect 15568 33847 15620 33856
rect 15568 33813 15577 33847
rect 15577 33813 15611 33847
rect 15611 33813 15620 33847
rect 15568 33804 15620 33813
rect 16580 33804 16632 33856
rect 16856 33847 16908 33856
rect 16856 33813 16865 33847
rect 16865 33813 16899 33847
rect 16899 33813 16908 33847
rect 16856 33804 16908 33813
rect 17592 33847 17644 33856
rect 17592 33813 17601 33847
rect 17601 33813 17635 33847
rect 17635 33813 17644 33847
rect 17592 33804 17644 33813
rect 18880 33847 18932 33856
rect 18880 33813 18889 33847
rect 18889 33813 18923 33847
rect 18923 33813 18932 33847
rect 18880 33804 18932 33813
rect 19800 33804 19852 33856
rect 22284 33847 22336 33856
rect 22284 33813 22293 33847
rect 22293 33813 22327 33847
rect 22327 33813 22336 33847
rect 22284 33804 22336 33813
rect 22836 33847 22888 33856
rect 22836 33813 22845 33847
rect 22845 33813 22879 33847
rect 22879 33813 22888 33847
rect 22836 33804 22888 33813
rect 23848 33804 23900 33856
rect 28540 33804 28592 33856
rect 29920 33804 29972 33856
rect 30104 33804 30156 33856
rect 32404 33872 32456 33924
rect 33048 33804 33100 33856
rect 4874 33702 4926 33754
rect 4938 33702 4990 33754
rect 5002 33702 5054 33754
rect 5066 33702 5118 33754
rect 5130 33702 5182 33754
rect 35594 33702 35646 33754
rect 35658 33702 35710 33754
rect 35722 33702 35774 33754
rect 35786 33702 35838 33754
rect 35850 33702 35902 33754
rect 9588 33643 9640 33652
rect 9588 33609 9597 33643
rect 9597 33609 9631 33643
rect 9631 33609 9640 33643
rect 9588 33600 9640 33609
rect 10508 33600 10560 33652
rect 6920 33532 6972 33584
rect 7380 33507 7432 33516
rect 7380 33473 7389 33507
rect 7389 33473 7423 33507
rect 7423 33473 7432 33507
rect 7380 33464 7432 33473
rect 8208 33532 8260 33584
rect 8392 33532 8444 33584
rect 10140 33532 10192 33584
rect 11796 33532 11848 33584
rect 12992 33532 13044 33584
rect 10048 33464 10100 33516
rect 16580 33600 16632 33652
rect 17500 33600 17552 33652
rect 18420 33600 18472 33652
rect 19064 33643 19116 33652
rect 19064 33609 19073 33643
rect 19073 33609 19107 33643
rect 19107 33609 19116 33643
rect 19064 33600 19116 33609
rect 22100 33600 22152 33652
rect 30104 33600 30156 33652
rect 32404 33643 32456 33652
rect 17592 33575 17644 33584
rect 17592 33541 17601 33575
rect 17601 33541 17635 33575
rect 17635 33541 17644 33575
rect 17592 33532 17644 33541
rect 17868 33532 17920 33584
rect 19432 33532 19484 33584
rect 17132 33464 17184 33516
rect 20720 33464 20772 33516
rect 21824 33464 21876 33516
rect 22284 33532 22336 33584
rect 24216 33507 24268 33516
rect 24216 33473 24225 33507
rect 24225 33473 24259 33507
rect 24259 33473 24268 33507
rect 24216 33464 24268 33473
rect 24860 33507 24912 33516
rect 24860 33473 24869 33507
rect 24869 33473 24903 33507
rect 24903 33473 24912 33507
rect 24860 33464 24912 33473
rect 26240 33464 26292 33516
rect 30012 33464 30064 33516
rect 32404 33609 32413 33643
rect 32413 33609 32447 33643
rect 32447 33609 32456 33643
rect 32404 33600 32456 33609
rect 33048 33643 33100 33652
rect 33048 33609 33057 33643
rect 33057 33609 33091 33643
rect 33091 33609 33100 33643
rect 33048 33600 33100 33609
rect 31392 33507 31444 33516
rect 8116 33439 8168 33448
rect 8116 33405 8125 33439
rect 8125 33405 8159 33439
rect 8159 33405 8168 33439
rect 8116 33396 8168 33405
rect 10968 33396 11020 33448
rect 12256 33439 12308 33448
rect 7012 33260 7064 33312
rect 12256 33405 12265 33439
rect 12265 33405 12299 33439
rect 12299 33405 12308 33439
rect 12256 33396 12308 33405
rect 12900 33396 12952 33448
rect 16028 33439 16080 33448
rect 16028 33405 16037 33439
rect 16037 33405 16071 33439
rect 16071 33405 16080 33439
rect 16028 33396 16080 33405
rect 16212 33439 16264 33448
rect 16212 33405 16221 33439
rect 16221 33405 16255 33439
rect 16255 33405 16264 33439
rect 16212 33396 16264 33405
rect 16672 33396 16724 33448
rect 22284 33439 22336 33448
rect 22284 33405 22293 33439
rect 22293 33405 22327 33439
rect 22327 33405 22336 33439
rect 22284 33396 22336 33405
rect 27712 33396 27764 33448
rect 26700 33328 26752 33380
rect 29000 33371 29052 33380
rect 29000 33337 29009 33371
rect 29009 33337 29043 33371
rect 29043 33337 29052 33371
rect 29000 33328 29052 33337
rect 29184 33439 29236 33448
rect 29184 33405 29193 33439
rect 29193 33405 29227 33439
rect 29227 33405 29236 33439
rect 29184 33396 29236 33405
rect 29920 33396 29972 33448
rect 31392 33473 31401 33507
rect 31401 33473 31435 33507
rect 31435 33473 31444 33507
rect 31392 33464 31444 33473
rect 29644 33328 29696 33380
rect 30380 33328 30432 33380
rect 33508 33464 33560 33516
rect 33784 33464 33836 33516
rect 14188 33260 14240 33312
rect 15108 33303 15160 33312
rect 15108 33269 15117 33303
rect 15117 33269 15151 33303
rect 15151 33269 15160 33303
rect 15108 33260 15160 33269
rect 23848 33260 23900 33312
rect 24952 33260 25004 33312
rect 27528 33260 27580 33312
rect 29184 33303 29236 33312
rect 29184 33269 29193 33303
rect 29193 33269 29227 33303
rect 29227 33269 29236 33303
rect 29184 33260 29236 33269
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 8484 33099 8536 33108
rect 8484 33065 8493 33099
rect 8493 33065 8527 33099
rect 8527 33065 8536 33099
rect 8484 33056 8536 33065
rect 9496 33056 9548 33108
rect 12072 33056 12124 33108
rect 14280 33056 14332 33108
rect 15108 33056 15160 33108
rect 17408 33056 17460 33108
rect 7012 32963 7064 32972
rect 7012 32929 7021 32963
rect 7021 32929 7055 32963
rect 7055 32929 7064 32963
rect 7012 32920 7064 32929
rect 10048 32963 10100 32972
rect 10048 32929 10057 32963
rect 10057 32929 10091 32963
rect 10091 32929 10100 32963
rect 10048 32920 10100 32929
rect 6460 32852 6512 32904
rect 6736 32895 6788 32904
rect 6736 32861 6745 32895
rect 6745 32861 6779 32895
rect 6779 32861 6788 32895
rect 6736 32852 6788 32861
rect 9680 32852 9732 32904
rect 10324 32920 10376 32972
rect 12624 32988 12676 33040
rect 12900 32920 12952 32972
rect 15568 32988 15620 33040
rect 11244 32852 11296 32904
rect 12348 32852 12400 32904
rect 12440 32852 12492 32904
rect 15200 32963 15252 32972
rect 15200 32929 15209 32963
rect 15209 32929 15243 32963
rect 15243 32929 15252 32963
rect 15200 32920 15252 32929
rect 16672 32920 16724 32972
rect 18420 32920 18472 32972
rect 19524 33056 19576 33108
rect 19800 33056 19852 33108
rect 24216 33056 24268 33108
rect 26240 33056 26292 33108
rect 26608 33056 26660 33108
rect 30104 33056 30156 33108
rect 30380 33056 30432 33108
rect 34520 33056 34572 33108
rect 27712 33031 27764 33040
rect 17960 32852 18012 32904
rect 22100 32920 22152 32972
rect 23940 32920 23992 32972
rect 25136 32963 25188 32972
rect 25136 32929 25145 32963
rect 25145 32929 25179 32963
rect 25179 32929 25188 32963
rect 25136 32920 25188 32929
rect 26700 32920 26752 32972
rect 21824 32895 21876 32904
rect 21824 32861 21833 32895
rect 21833 32861 21867 32895
rect 21867 32861 21876 32895
rect 21824 32852 21876 32861
rect 23848 32852 23900 32904
rect 26608 32852 26660 32904
rect 7288 32784 7340 32836
rect 12164 32784 12216 32836
rect 16856 32784 16908 32836
rect 18880 32784 18932 32836
rect 20444 32784 20496 32836
rect 25320 32784 25372 32836
rect 27712 32997 27721 33031
rect 27721 32997 27755 33031
rect 27755 32997 27764 33031
rect 27712 32988 27764 32997
rect 30012 32988 30064 33040
rect 28356 32920 28408 32972
rect 29184 32920 29236 32972
rect 31300 32988 31352 33040
rect 31392 32988 31444 33040
rect 27988 32852 28040 32904
rect 28632 32895 28684 32904
rect 28632 32861 28641 32895
rect 28641 32861 28675 32895
rect 28675 32861 28684 32895
rect 28632 32852 28684 32861
rect 29368 32852 29420 32904
rect 33508 32920 33560 32972
rect 32772 32895 32824 32904
rect 32772 32861 32781 32895
rect 32781 32861 32815 32895
rect 32815 32861 32824 32895
rect 32772 32852 32824 32861
rect 11060 32759 11112 32768
rect 11060 32725 11069 32759
rect 11069 32725 11103 32759
rect 11103 32725 11112 32759
rect 11060 32716 11112 32725
rect 11520 32716 11572 32768
rect 13360 32716 13412 32768
rect 15200 32716 15252 32768
rect 16028 32716 16080 32768
rect 17500 32716 17552 32768
rect 17868 32716 17920 32768
rect 18512 32759 18564 32768
rect 18512 32725 18521 32759
rect 18521 32725 18555 32759
rect 18555 32725 18564 32759
rect 18512 32716 18564 32725
rect 23204 32759 23256 32768
rect 23204 32725 23213 32759
rect 23213 32725 23247 32759
rect 23247 32725 23256 32759
rect 23204 32716 23256 32725
rect 24952 32759 25004 32768
rect 24952 32725 24961 32759
rect 24961 32725 24995 32759
rect 24995 32725 25004 32759
rect 24952 32716 25004 32725
rect 28264 32716 28316 32768
rect 32036 32784 32088 32836
rect 33048 32784 33100 32836
rect 33140 32784 33192 32836
rect 4874 32614 4926 32666
rect 4938 32614 4990 32666
rect 5002 32614 5054 32666
rect 5066 32614 5118 32666
rect 5130 32614 5182 32666
rect 35594 32614 35646 32666
rect 35658 32614 35710 32666
rect 35722 32614 35774 32666
rect 35786 32614 35838 32666
rect 35850 32614 35902 32666
rect 8116 32512 8168 32564
rect 8300 32444 8352 32496
rect 7840 32308 7892 32360
rect 9404 32512 9456 32564
rect 15200 32512 15252 32564
rect 18512 32512 18564 32564
rect 19800 32512 19852 32564
rect 20444 32555 20496 32564
rect 20444 32521 20453 32555
rect 20453 32521 20487 32555
rect 20487 32521 20496 32555
rect 20444 32512 20496 32521
rect 22284 32512 22336 32564
rect 23388 32512 23440 32564
rect 11060 32444 11112 32496
rect 8944 32376 8996 32428
rect 9312 32419 9364 32428
rect 9312 32385 9321 32419
rect 9321 32385 9355 32419
rect 9355 32385 9364 32419
rect 9312 32376 9364 32385
rect 10968 32419 11020 32428
rect 10968 32385 10977 32419
rect 10977 32385 11011 32419
rect 11011 32385 11020 32419
rect 10968 32376 11020 32385
rect 12072 32419 12124 32428
rect 12072 32385 12081 32419
rect 12081 32385 12115 32419
rect 12115 32385 12124 32419
rect 12072 32376 12124 32385
rect 12348 32376 12400 32428
rect 16856 32376 16908 32428
rect 18052 32419 18104 32428
rect 18052 32385 18061 32419
rect 18061 32385 18095 32419
rect 18095 32385 18104 32419
rect 18052 32376 18104 32385
rect 19524 32419 19576 32428
rect 19524 32385 19533 32419
rect 19533 32385 19567 32419
rect 19567 32385 19576 32419
rect 19524 32376 19576 32385
rect 21272 32419 21324 32428
rect 9128 32308 9180 32360
rect 12164 32351 12216 32360
rect 12164 32317 12173 32351
rect 12173 32317 12207 32351
rect 12207 32317 12216 32351
rect 12164 32308 12216 32317
rect 12624 32308 12676 32360
rect 15200 32308 15252 32360
rect 16672 32308 16724 32360
rect 17132 32308 17184 32360
rect 19708 32351 19760 32360
rect 19708 32317 19717 32351
rect 19717 32317 19751 32351
rect 19751 32317 19760 32351
rect 19708 32308 19760 32317
rect 20076 32308 20128 32360
rect 21272 32385 21281 32419
rect 21281 32385 21315 32419
rect 21315 32385 21324 32419
rect 21272 32376 21324 32385
rect 22192 32419 22244 32428
rect 22192 32385 22201 32419
rect 22201 32385 22235 32419
rect 22235 32385 22244 32419
rect 22192 32376 22244 32385
rect 22836 32419 22888 32428
rect 22836 32385 22845 32419
rect 22845 32385 22879 32419
rect 22879 32385 22888 32419
rect 22836 32376 22888 32385
rect 20904 32308 20956 32360
rect 22284 32308 22336 32360
rect 23940 32351 23992 32360
rect 12348 32240 12400 32292
rect 23940 32317 23949 32351
rect 23949 32317 23983 32351
rect 23983 32317 23992 32351
rect 23940 32308 23992 32317
rect 25136 32444 25188 32496
rect 29000 32512 29052 32564
rect 29552 32512 29604 32564
rect 30932 32512 30984 32564
rect 33048 32555 33100 32564
rect 33048 32521 33057 32555
rect 33057 32521 33091 32555
rect 33091 32521 33100 32555
rect 33048 32512 33100 32521
rect 27528 32444 27580 32496
rect 29644 32487 29696 32496
rect 26608 32376 26660 32428
rect 27712 32376 27764 32428
rect 25320 32308 25372 32360
rect 25044 32240 25096 32292
rect 6644 32172 6696 32224
rect 8668 32215 8720 32224
rect 8668 32181 8677 32215
rect 8677 32181 8711 32215
rect 8711 32181 8720 32215
rect 8668 32172 8720 32181
rect 9220 32215 9272 32224
rect 9220 32181 9229 32215
rect 9229 32181 9263 32215
rect 9263 32181 9272 32215
rect 9220 32172 9272 32181
rect 10508 32172 10560 32224
rect 11152 32215 11204 32224
rect 11152 32181 11161 32215
rect 11161 32181 11195 32215
rect 11195 32181 11204 32215
rect 11152 32172 11204 32181
rect 11704 32215 11756 32224
rect 11704 32181 11713 32215
rect 11713 32181 11747 32215
rect 11747 32181 11756 32215
rect 11704 32172 11756 32181
rect 14464 32172 14516 32224
rect 17316 32172 17368 32224
rect 18512 32172 18564 32224
rect 21456 32172 21508 32224
rect 22008 32215 22060 32224
rect 22008 32181 22017 32215
rect 22017 32181 22051 32215
rect 22051 32181 22060 32215
rect 22008 32172 22060 32181
rect 23296 32215 23348 32224
rect 23296 32181 23305 32215
rect 23305 32181 23339 32215
rect 23339 32181 23348 32215
rect 23296 32172 23348 32181
rect 24952 32172 25004 32224
rect 26424 32215 26476 32224
rect 26424 32181 26433 32215
rect 26433 32181 26467 32215
rect 26467 32181 26476 32215
rect 26424 32172 26476 32181
rect 27712 32172 27764 32224
rect 29644 32453 29653 32487
rect 29653 32453 29687 32487
rect 29687 32453 29696 32487
rect 29644 32444 29696 32453
rect 29920 32419 29972 32428
rect 29920 32385 29929 32419
rect 29929 32385 29963 32419
rect 29963 32385 29972 32419
rect 29920 32376 29972 32385
rect 31116 32419 31168 32428
rect 31116 32385 31125 32419
rect 31125 32385 31159 32419
rect 31159 32385 31168 32419
rect 31116 32376 31168 32385
rect 31300 32376 31352 32428
rect 32036 32444 32088 32496
rect 33784 32419 33836 32428
rect 31300 32240 31352 32292
rect 32404 32283 32456 32292
rect 32404 32249 32413 32283
rect 32413 32249 32447 32283
rect 32447 32249 32456 32283
rect 32404 32240 32456 32249
rect 30012 32172 30064 32224
rect 30840 32172 30892 32224
rect 31484 32172 31536 32224
rect 33784 32385 33793 32419
rect 33793 32385 33827 32419
rect 33827 32385 33836 32419
rect 33784 32376 33836 32385
rect 33692 32215 33744 32224
rect 33692 32181 33701 32215
rect 33701 32181 33735 32215
rect 33735 32181 33744 32215
rect 33692 32172 33744 32181
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 7288 32011 7340 32020
rect 7288 31977 7297 32011
rect 7297 31977 7331 32011
rect 7331 31977 7340 32011
rect 7288 31968 7340 31977
rect 7840 32011 7892 32020
rect 7840 31977 7849 32011
rect 7849 31977 7883 32011
rect 7883 31977 7892 32011
rect 7840 31968 7892 31977
rect 11060 31968 11112 32020
rect 11152 31968 11204 32020
rect 12348 31968 12400 32020
rect 15016 32011 15068 32020
rect 11520 31943 11572 31952
rect 11520 31909 11529 31943
rect 11529 31909 11563 31943
rect 11563 31909 11572 31943
rect 11520 31900 11572 31909
rect 15016 31977 15025 32011
rect 15025 31977 15059 32011
rect 15059 31977 15068 32011
rect 15016 31968 15068 31977
rect 22008 31968 22060 32020
rect 22192 31968 22244 32020
rect 29276 31968 29328 32020
rect 30932 31968 30984 32020
rect 8024 31832 8076 31884
rect 8668 31832 8720 31884
rect 12256 31832 12308 31884
rect 14280 31832 14332 31884
rect 22100 31900 22152 31952
rect 23388 31900 23440 31952
rect 16120 31875 16172 31884
rect 16120 31841 16129 31875
rect 16129 31841 16163 31875
rect 16163 31841 16172 31875
rect 16120 31832 16172 31841
rect 19524 31832 19576 31884
rect 19892 31832 19944 31884
rect 22560 31832 22612 31884
rect 24952 31875 25004 31884
rect 24952 31841 24961 31875
rect 24961 31841 24995 31875
rect 24995 31841 25004 31875
rect 24952 31832 25004 31841
rect 25320 31832 25372 31884
rect 27896 31832 27948 31884
rect 1952 31764 2004 31816
rect 6920 31764 6972 31816
rect 7104 31764 7156 31816
rect 9128 31807 9180 31816
rect 9128 31773 9137 31807
rect 9137 31773 9171 31807
rect 9171 31773 9180 31807
rect 9128 31764 9180 31773
rect 9772 31807 9824 31816
rect 9772 31773 9781 31807
rect 9781 31773 9815 31807
rect 9815 31773 9824 31807
rect 9772 31764 9824 31773
rect 13360 31764 13412 31816
rect 10508 31696 10560 31748
rect 16028 31764 16080 31816
rect 17132 31807 17184 31816
rect 17132 31773 17141 31807
rect 17141 31773 17175 31807
rect 17175 31773 17184 31807
rect 17132 31764 17184 31773
rect 18512 31764 18564 31816
rect 19616 31807 19668 31816
rect 19616 31773 19625 31807
rect 19625 31773 19659 31807
rect 19659 31773 19668 31807
rect 19616 31764 19668 31773
rect 20076 31807 20128 31816
rect 20076 31773 20085 31807
rect 20085 31773 20119 31807
rect 20119 31773 20128 31807
rect 20076 31764 20128 31773
rect 20352 31764 20404 31816
rect 23204 31764 23256 31816
rect 23388 31807 23440 31816
rect 23388 31773 23397 31807
rect 23397 31773 23431 31807
rect 23431 31773 23440 31807
rect 24676 31807 24728 31816
rect 23388 31764 23440 31773
rect 24676 31773 24685 31807
rect 24685 31773 24719 31807
rect 24719 31773 24728 31807
rect 24676 31764 24728 31773
rect 27620 31807 27672 31816
rect 1584 31671 1636 31680
rect 1584 31637 1593 31671
rect 1593 31637 1627 31671
rect 1627 31637 1636 31671
rect 1584 31628 1636 31637
rect 6552 31628 6604 31680
rect 8208 31671 8260 31680
rect 8208 31637 8217 31671
rect 8217 31637 8251 31671
rect 8251 31637 8260 31671
rect 8208 31628 8260 31637
rect 8300 31671 8352 31680
rect 8300 31637 8309 31671
rect 8309 31637 8343 31671
rect 8343 31637 8352 31671
rect 8300 31628 8352 31637
rect 14004 31628 14056 31680
rect 15568 31671 15620 31680
rect 15568 31637 15577 31671
rect 15577 31637 15611 31671
rect 15611 31637 15620 31671
rect 15568 31628 15620 31637
rect 16028 31671 16080 31680
rect 16028 31637 16037 31671
rect 16037 31637 16071 31671
rect 16071 31637 16080 31671
rect 16028 31628 16080 31637
rect 17408 31739 17460 31748
rect 17408 31705 17417 31739
rect 17417 31705 17451 31739
rect 17451 31705 17460 31739
rect 17408 31696 17460 31705
rect 17684 31628 17736 31680
rect 17776 31628 17828 31680
rect 19432 31671 19484 31680
rect 19432 31637 19441 31671
rect 19441 31637 19475 31671
rect 19475 31637 19484 31671
rect 19432 31628 19484 31637
rect 21456 31696 21508 31748
rect 26608 31696 26660 31748
rect 27620 31773 27629 31807
rect 27629 31773 27663 31807
rect 27663 31773 27672 31807
rect 27620 31764 27672 31773
rect 28080 31807 28132 31816
rect 28080 31773 28089 31807
rect 28089 31773 28123 31807
rect 28123 31773 28132 31807
rect 28080 31764 28132 31773
rect 28632 31764 28684 31816
rect 29092 31900 29144 31952
rect 29368 31900 29420 31952
rect 28172 31696 28224 31748
rect 29000 31764 29052 31816
rect 29552 31764 29604 31816
rect 30748 31832 30800 31884
rect 32772 31832 32824 31884
rect 33324 31832 33376 31884
rect 30656 31764 30708 31816
rect 30932 31764 30984 31816
rect 33784 31807 33836 31816
rect 33784 31773 33793 31807
rect 33793 31773 33827 31807
rect 33827 31773 33836 31807
rect 33784 31764 33836 31773
rect 34520 31764 34572 31816
rect 31576 31739 31628 31748
rect 26884 31628 26936 31680
rect 29736 31628 29788 31680
rect 29920 31628 29972 31680
rect 31576 31705 31585 31739
rect 31585 31705 31619 31739
rect 31619 31705 31628 31739
rect 31576 31696 31628 31705
rect 32404 31628 32456 31680
rect 37096 31671 37148 31680
rect 37096 31637 37105 31671
rect 37105 31637 37139 31671
rect 37139 31637 37148 31671
rect 37096 31628 37148 31637
rect 4874 31526 4926 31578
rect 4938 31526 4990 31578
rect 5002 31526 5054 31578
rect 5066 31526 5118 31578
rect 5130 31526 5182 31578
rect 35594 31526 35646 31578
rect 35658 31526 35710 31578
rect 35722 31526 35774 31578
rect 35786 31526 35838 31578
rect 35850 31526 35902 31578
rect 8944 31424 8996 31476
rect 11704 31424 11756 31476
rect 9220 31356 9272 31408
rect 11520 31356 11572 31408
rect 17408 31424 17460 31476
rect 19064 31467 19116 31476
rect 19064 31433 19073 31467
rect 19073 31433 19107 31467
rect 19107 31433 19116 31467
rect 19064 31424 19116 31433
rect 23296 31424 23348 31476
rect 15292 31356 15344 31408
rect 16028 31356 16080 31408
rect 17224 31356 17276 31408
rect 17776 31356 17828 31408
rect 25044 31424 25096 31476
rect 7012 31331 7064 31340
rect 7012 31297 7021 31331
rect 7021 31297 7055 31331
rect 7055 31297 7064 31331
rect 7012 31288 7064 31297
rect 11888 31288 11940 31340
rect 11980 31288 12032 31340
rect 6460 31220 6512 31272
rect 10876 31220 10928 31272
rect 12256 31220 12308 31272
rect 13820 31220 13872 31272
rect 17868 31288 17920 31340
rect 19892 31288 19944 31340
rect 20904 31288 20956 31340
rect 21272 31331 21324 31340
rect 21272 31297 21281 31331
rect 21281 31297 21315 31331
rect 21315 31297 21324 31331
rect 21272 31288 21324 31297
rect 19156 31263 19208 31272
rect 19156 31229 19165 31263
rect 19165 31229 19199 31263
rect 19199 31229 19208 31263
rect 19156 31220 19208 31229
rect 19340 31263 19392 31272
rect 19340 31229 19349 31263
rect 19349 31229 19383 31263
rect 19383 31229 19392 31263
rect 19340 31220 19392 31229
rect 9404 31127 9456 31136
rect 9404 31093 9413 31127
rect 9413 31093 9447 31127
rect 9447 31093 9456 31127
rect 9404 31084 9456 31093
rect 16580 31084 16632 31136
rect 17960 31084 18012 31136
rect 26424 31356 26476 31408
rect 23848 31288 23900 31340
rect 24584 31288 24636 31340
rect 22652 31263 22704 31272
rect 22652 31229 22661 31263
rect 22661 31229 22695 31263
rect 22695 31229 22704 31263
rect 22652 31220 22704 31229
rect 22928 31220 22980 31272
rect 24676 31263 24728 31272
rect 24676 31229 24685 31263
rect 24685 31229 24719 31263
rect 24719 31229 24728 31263
rect 24676 31220 24728 31229
rect 21364 31127 21416 31136
rect 21364 31093 21373 31127
rect 21373 31093 21407 31127
rect 21407 31093 21416 31127
rect 21364 31084 21416 31093
rect 23572 31084 23624 31136
rect 29000 31424 29052 31476
rect 26884 31356 26936 31408
rect 33600 31424 33652 31476
rect 34520 31424 34572 31476
rect 36912 31424 36964 31476
rect 27988 31331 28040 31340
rect 27988 31297 27997 31331
rect 27997 31297 28031 31331
rect 28031 31297 28040 31331
rect 27988 31288 28040 31297
rect 31116 31356 31168 31408
rect 31300 31356 31352 31408
rect 31484 31356 31536 31408
rect 31668 31356 31720 31408
rect 27620 31152 27672 31204
rect 29276 31152 29328 31204
rect 30840 31195 30892 31204
rect 30840 31161 30849 31195
rect 30849 31161 30883 31195
rect 30883 31161 30892 31195
rect 30840 31152 30892 31161
rect 27896 31127 27948 31136
rect 27896 31093 27905 31127
rect 27905 31093 27939 31127
rect 27939 31093 27948 31127
rect 27896 31084 27948 31093
rect 28448 31084 28500 31136
rect 30748 31084 30800 31136
rect 30932 31084 30984 31136
rect 34336 31288 34388 31340
rect 33600 31084 33652 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 8208 30923 8260 30932
rect 8208 30889 8217 30923
rect 8217 30889 8251 30923
rect 8251 30889 8260 30923
rect 8208 30880 8260 30889
rect 10968 30880 11020 30932
rect 11888 30880 11940 30932
rect 16028 30880 16080 30932
rect 16120 30880 16172 30932
rect 19340 30880 19392 30932
rect 19616 30880 19668 30932
rect 23848 30880 23900 30932
rect 24584 30923 24636 30932
rect 24584 30889 24593 30923
rect 24593 30889 24627 30923
rect 24627 30889 24636 30923
rect 24584 30880 24636 30889
rect 27988 30880 28040 30932
rect 29736 30923 29788 30932
rect 12624 30812 12676 30864
rect 15108 30812 15160 30864
rect 7104 30744 7156 30796
rect 9772 30744 9824 30796
rect 11520 30744 11572 30796
rect 12532 30744 12584 30796
rect 14832 30744 14884 30796
rect 17316 30744 17368 30796
rect 21272 30812 21324 30864
rect 28080 30812 28132 30864
rect 28908 30855 28960 30864
rect 28908 30821 28917 30855
rect 28917 30821 28951 30855
rect 28951 30821 28960 30855
rect 28908 30812 28960 30821
rect 29736 30889 29745 30923
rect 29745 30889 29779 30923
rect 29779 30889 29788 30923
rect 29736 30880 29788 30889
rect 30564 30880 30616 30932
rect 31208 30880 31260 30932
rect 34336 30923 34388 30932
rect 34336 30889 34345 30923
rect 34345 30889 34379 30923
rect 34379 30889 34388 30923
rect 34336 30880 34388 30889
rect 30840 30812 30892 30864
rect 19892 30787 19944 30796
rect 19892 30753 19901 30787
rect 19901 30753 19935 30787
rect 19935 30753 19944 30787
rect 19892 30744 19944 30753
rect 19984 30787 20036 30796
rect 19984 30753 19993 30787
rect 19993 30753 20027 30787
rect 20027 30753 20036 30787
rect 19984 30744 20036 30753
rect 22192 30744 22244 30796
rect 24860 30744 24912 30796
rect 25136 30787 25188 30796
rect 25136 30753 25145 30787
rect 25145 30753 25179 30787
rect 25179 30753 25188 30787
rect 25136 30744 25188 30753
rect 29920 30744 29972 30796
rect 30748 30744 30800 30796
rect 32404 30744 32456 30796
rect 33600 30744 33652 30796
rect 6460 30719 6512 30728
rect 6460 30685 6469 30719
rect 6469 30685 6503 30719
rect 6503 30685 6512 30719
rect 6460 30676 6512 30685
rect 9220 30719 9272 30728
rect 9220 30685 9229 30719
rect 9229 30685 9263 30719
rect 9263 30685 9272 30719
rect 9220 30676 9272 30685
rect 12164 30719 12216 30728
rect 12164 30685 12173 30719
rect 12173 30685 12207 30719
rect 12207 30685 12216 30719
rect 12164 30676 12216 30685
rect 15568 30676 15620 30728
rect 17684 30719 17736 30728
rect 17684 30685 17693 30719
rect 17693 30685 17727 30719
rect 17727 30685 17736 30719
rect 17684 30676 17736 30685
rect 18512 30676 18564 30728
rect 19156 30676 19208 30728
rect 20812 30676 20864 30728
rect 22928 30719 22980 30728
rect 22928 30685 22937 30719
rect 22937 30685 22971 30719
rect 22971 30685 22980 30719
rect 23572 30719 23624 30728
rect 22928 30676 22980 30685
rect 23572 30685 23581 30719
rect 23581 30685 23615 30719
rect 23615 30685 23624 30719
rect 23572 30676 23624 30685
rect 24952 30719 25004 30728
rect 24952 30685 24961 30719
rect 24961 30685 24995 30719
rect 24995 30685 25004 30719
rect 24952 30676 25004 30685
rect 25964 30719 26016 30728
rect 25964 30685 25973 30719
rect 25973 30685 26007 30719
rect 26007 30685 26016 30719
rect 25964 30676 26016 30685
rect 26608 30719 26660 30728
rect 26608 30685 26617 30719
rect 26617 30685 26651 30719
rect 26651 30685 26660 30719
rect 26608 30676 26660 30685
rect 27344 30719 27396 30728
rect 27344 30685 27353 30719
rect 27353 30685 27387 30719
rect 27387 30685 27396 30719
rect 27344 30676 27396 30685
rect 6644 30608 6696 30660
rect 6552 30540 6604 30592
rect 11980 30608 12032 30660
rect 13636 30651 13688 30660
rect 13636 30617 13645 30651
rect 13645 30617 13679 30651
rect 13679 30617 13688 30651
rect 13636 30608 13688 30617
rect 9312 30583 9364 30592
rect 9312 30549 9321 30583
rect 9321 30549 9355 30583
rect 9355 30549 9364 30583
rect 9312 30540 9364 30549
rect 16396 30608 16448 30660
rect 21364 30608 21416 30660
rect 16580 30540 16632 30592
rect 23848 30608 23900 30660
rect 27252 30608 27304 30660
rect 27620 30719 27672 30728
rect 27620 30685 27629 30719
rect 27629 30685 27663 30719
rect 27663 30685 27672 30719
rect 27620 30676 27672 30685
rect 27896 30676 27948 30728
rect 27988 30676 28040 30728
rect 28448 30719 28500 30728
rect 28448 30685 28457 30719
rect 28457 30685 28491 30719
rect 28491 30685 28500 30719
rect 28448 30676 28500 30685
rect 29000 30676 29052 30728
rect 33692 30608 33744 30660
rect 25228 30540 25280 30592
rect 26516 30583 26568 30592
rect 26516 30549 26525 30583
rect 26525 30549 26559 30583
rect 26559 30549 26568 30583
rect 26516 30540 26568 30549
rect 27804 30540 27856 30592
rect 28448 30540 28500 30592
rect 33968 30583 34020 30592
rect 33968 30549 33977 30583
rect 33977 30549 34011 30583
rect 34011 30549 34020 30583
rect 33968 30540 34020 30549
rect 4874 30438 4926 30490
rect 4938 30438 4990 30490
rect 5002 30438 5054 30490
rect 5066 30438 5118 30490
rect 5130 30438 5182 30490
rect 35594 30438 35646 30490
rect 35658 30438 35710 30490
rect 35722 30438 35774 30490
rect 35786 30438 35838 30490
rect 35850 30438 35902 30490
rect 8300 30336 8352 30388
rect 9404 30336 9456 30388
rect 11152 30336 11204 30388
rect 12532 30336 12584 30388
rect 16580 30336 16632 30388
rect 8208 30268 8260 30320
rect 12900 30268 12952 30320
rect 14832 30311 14884 30320
rect 14832 30277 14841 30311
rect 14841 30277 14875 30311
rect 14875 30277 14884 30311
rect 14832 30268 14884 30277
rect 16396 30268 16448 30320
rect 17224 30311 17276 30320
rect 17224 30277 17233 30311
rect 17233 30277 17267 30311
rect 17267 30277 17276 30311
rect 17224 30268 17276 30277
rect 19064 30336 19116 30388
rect 17684 30268 17736 30320
rect 7012 30064 7064 30116
rect 8300 30200 8352 30252
rect 11244 30200 11296 30252
rect 12072 30200 12124 30252
rect 8208 30132 8260 30184
rect 9588 30132 9640 30184
rect 11152 30132 11204 30184
rect 12256 30132 12308 30184
rect 9128 30064 9180 30116
rect 12992 30200 13044 30252
rect 14924 30200 14976 30252
rect 15108 30200 15160 30252
rect 15752 30200 15804 30252
rect 17040 30200 17092 30252
rect 18052 30200 18104 30252
rect 18512 30243 18564 30252
rect 18512 30209 18521 30243
rect 18521 30209 18555 30243
rect 18555 30209 18564 30243
rect 18512 30200 18564 30209
rect 19432 30268 19484 30320
rect 20352 30268 20404 30320
rect 20812 30268 20864 30320
rect 22284 30268 22336 30320
rect 25964 30336 26016 30388
rect 27344 30336 27396 30388
rect 28356 30336 28408 30388
rect 28448 30268 28500 30320
rect 28908 30336 28960 30388
rect 29276 30336 29328 30388
rect 22376 30200 22428 30252
rect 23848 30243 23900 30252
rect 12440 30132 12492 30184
rect 14280 30132 14332 30184
rect 15568 30132 15620 30184
rect 16212 30132 16264 30184
rect 19984 30132 20036 30184
rect 20812 30175 20864 30184
rect 20812 30141 20821 30175
rect 20821 30141 20855 30175
rect 20855 30141 20864 30175
rect 20812 30132 20864 30141
rect 23848 30209 23857 30243
rect 23857 30209 23891 30243
rect 23891 30209 23900 30243
rect 23848 30200 23900 30209
rect 25044 30243 25096 30252
rect 25044 30209 25053 30243
rect 25053 30209 25087 30243
rect 25087 30209 25096 30243
rect 25044 30200 25096 30209
rect 26792 30200 26844 30252
rect 27252 30200 27304 30252
rect 23756 30132 23808 30184
rect 24032 30175 24084 30184
rect 24032 30141 24041 30175
rect 24041 30141 24075 30175
rect 24075 30141 24084 30175
rect 24032 30132 24084 30141
rect 24860 30175 24912 30184
rect 24860 30141 24869 30175
rect 24869 30141 24903 30175
rect 24903 30141 24912 30175
rect 24860 30132 24912 30141
rect 10140 29996 10192 30048
rect 11612 29996 11664 30048
rect 15292 30039 15344 30048
rect 15292 30005 15301 30039
rect 15301 30005 15335 30039
rect 15335 30005 15344 30039
rect 15292 29996 15344 30005
rect 16856 30039 16908 30048
rect 16856 30005 16865 30039
rect 16865 30005 16899 30039
rect 16899 30005 16908 30039
rect 16856 29996 16908 30005
rect 23572 30064 23624 30116
rect 27620 30064 27672 30116
rect 21180 29996 21232 30048
rect 23480 30039 23532 30048
rect 23480 30005 23489 30039
rect 23489 30005 23523 30039
rect 23523 30005 23532 30039
rect 23480 29996 23532 30005
rect 24860 29996 24912 30048
rect 28172 30200 28224 30252
rect 28540 30243 28592 30252
rect 28540 30209 28544 30243
rect 28544 30209 28578 30243
rect 28578 30209 28592 30243
rect 28540 30200 28592 30209
rect 28632 30243 28684 30252
rect 28632 30209 28641 30243
rect 28641 30209 28675 30243
rect 28675 30209 28684 30243
rect 28632 30200 28684 30209
rect 28816 30243 28868 30252
rect 28816 30209 28861 30243
rect 28861 30209 28868 30243
rect 28816 30200 28868 30209
rect 30932 30200 30984 30252
rect 31484 30243 31536 30252
rect 31484 30209 31493 30243
rect 31493 30209 31527 30243
rect 31527 30209 31536 30243
rect 31484 30200 31536 30209
rect 32128 30200 32180 30252
rect 33048 30200 33100 30252
rect 33968 30200 34020 30252
rect 30564 30175 30616 30184
rect 30564 30141 30573 30175
rect 30573 30141 30607 30175
rect 30607 30141 30616 30175
rect 30564 30132 30616 30141
rect 31576 30132 31628 30184
rect 33324 30132 33376 30184
rect 27896 30064 27948 30116
rect 28080 29996 28132 30048
rect 28356 30039 28408 30048
rect 28356 30005 28365 30039
rect 28365 30005 28399 30039
rect 28399 30005 28408 30039
rect 28356 29996 28408 30005
rect 28908 30064 28960 30116
rect 29092 30064 29144 30116
rect 29736 29996 29788 30048
rect 34428 29996 34480 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 6920 29792 6972 29844
rect 8024 29724 8076 29776
rect 8300 29699 8352 29708
rect 8300 29665 8309 29699
rect 8309 29665 8343 29699
rect 8343 29665 8352 29699
rect 8300 29656 8352 29665
rect 6920 29588 6972 29640
rect 8760 29792 8812 29844
rect 9220 29792 9272 29844
rect 12900 29835 12952 29844
rect 11152 29724 11204 29776
rect 10876 29656 10928 29708
rect 11060 29656 11112 29708
rect 12900 29801 12909 29835
rect 12909 29801 12943 29835
rect 12943 29801 12952 29835
rect 12900 29792 12952 29801
rect 15568 29792 15620 29844
rect 15752 29835 15804 29844
rect 15752 29801 15761 29835
rect 15761 29801 15795 29835
rect 15795 29801 15804 29835
rect 15752 29792 15804 29801
rect 19708 29835 19760 29844
rect 13636 29724 13688 29776
rect 19708 29801 19717 29835
rect 19717 29801 19751 29835
rect 19751 29801 19760 29835
rect 19708 29792 19760 29801
rect 22284 29792 22336 29844
rect 22376 29792 22428 29844
rect 25044 29792 25096 29844
rect 27436 29792 27488 29844
rect 28908 29792 28960 29844
rect 6092 29495 6144 29504
rect 6092 29461 6101 29495
rect 6101 29461 6135 29495
rect 6135 29461 6144 29495
rect 6092 29452 6144 29461
rect 7288 29452 7340 29504
rect 8116 29452 8168 29504
rect 8392 29452 8444 29504
rect 10140 29631 10192 29640
rect 10140 29597 10149 29631
rect 10149 29597 10183 29631
rect 10183 29597 10192 29631
rect 10140 29588 10192 29597
rect 11152 29631 11204 29640
rect 11152 29597 11161 29631
rect 11161 29597 11195 29631
rect 11195 29597 11204 29631
rect 11152 29588 11204 29597
rect 18144 29656 18196 29708
rect 17500 29588 17552 29640
rect 18512 29588 18564 29640
rect 18604 29588 18656 29640
rect 27712 29724 27764 29776
rect 22928 29656 22980 29708
rect 23572 29699 23624 29708
rect 23572 29665 23581 29699
rect 23581 29665 23615 29699
rect 23615 29665 23624 29699
rect 23572 29656 23624 29665
rect 23664 29699 23716 29708
rect 23664 29665 23673 29699
rect 23673 29665 23707 29699
rect 23707 29665 23716 29699
rect 25228 29699 25280 29708
rect 23664 29656 23716 29665
rect 25228 29665 25237 29699
rect 25237 29665 25271 29699
rect 25271 29665 25280 29699
rect 25228 29656 25280 29665
rect 27988 29699 28040 29708
rect 27988 29665 27997 29699
rect 27997 29665 28031 29699
rect 28031 29665 28040 29699
rect 27988 29656 28040 29665
rect 28264 29724 28316 29776
rect 29920 29724 29972 29776
rect 33048 29835 33100 29844
rect 33048 29801 33057 29835
rect 33057 29801 33091 29835
rect 33091 29801 33100 29835
rect 33048 29792 33100 29801
rect 28448 29656 28500 29708
rect 29000 29656 29052 29708
rect 33968 29656 34020 29708
rect 14648 29563 14700 29572
rect 14648 29529 14657 29563
rect 14657 29529 14691 29563
rect 14691 29529 14700 29563
rect 14648 29520 14700 29529
rect 15476 29520 15528 29572
rect 19616 29520 19668 29572
rect 23480 29631 23532 29640
rect 23480 29597 23489 29631
rect 23489 29597 23523 29631
rect 23523 29597 23532 29631
rect 23480 29588 23532 29597
rect 24860 29588 24912 29640
rect 27804 29588 27856 29640
rect 27896 29631 27948 29640
rect 27896 29597 27905 29631
rect 27905 29597 27939 29631
rect 27939 29597 27948 29631
rect 27896 29588 27948 29597
rect 21180 29563 21232 29572
rect 13636 29495 13688 29504
rect 13636 29461 13645 29495
rect 13645 29461 13679 29495
rect 13679 29461 13688 29495
rect 13636 29452 13688 29461
rect 16120 29495 16172 29504
rect 16120 29461 16129 29495
rect 16129 29461 16163 29495
rect 16163 29461 16172 29495
rect 16120 29452 16172 29461
rect 16304 29452 16356 29504
rect 18420 29495 18472 29504
rect 18420 29461 18429 29495
rect 18429 29461 18463 29495
rect 18463 29461 18472 29495
rect 18420 29452 18472 29461
rect 18512 29495 18564 29504
rect 18512 29461 18521 29495
rect 18521 29461 18555 29495
rect 18555 29461 18564 29495
rect 18512 29452 18564 29461
rect 20260 29452 20312 29504
rect 21180 29529 21189 29563
rect 21189 29529 21223 29563
rect 21223 29529 21232 29563
rect 21180 29520 21232 29529
rect 21640 29520 21692 29572
rect 26516 29520 26568 29572
rect 28080 29520 28132 29572
rect 28816 29588 28868 29640
rect 29092 29631 29144 29640
rect 29092 29597 29101 29631
rect 29101 29597 29135 29631
rect 29135 29597 29144 29631
rect 29092 29588 29144 29597
rect 29184 29631 29236 29640
rect 29184 29597 29193 29631
rect 29193 29597 29227 29631
rect 29227 29597 29236 29631
rect 29184 29588 29236 29597
rect 29552 29588 29604 29640
rect 29828 29588 29880 29640
rect 32036 29588 32088 29640
rect 32220 29631 32272 29640
rect 32220 29597 32229 29631
rect 32229 29597 32263 29631
rect 32263 29597 32272 29631
rect 32220 29588 32272 29597
rect 30012 29563 30064 29572
rect 30012 29529 30021 29563
rect 30021 29529 30055 29563
rect 30055 29529 30064 29563
rect 30748 29563 30800 29572
rect 30012 29520 30064 29529
rect 30748 29529 30757 29563
rect 30757 29529 30791 29563
rect 30791 29529 30800 29563
rect 30748 29520 30800 29529
rect 33416 29520 33468 29572
rect 26792 29452 26844 29504
rect 29736 29452 29788 29504
rect 30656 29452 30708 29504
rect 31116 29495 31168 29504
rect 31116 29461 31125 29495
rect 31125 29461 31159 29495
rect 31159 29461 31168 29495
rect 31116 29452 31168 29461
rect 32404 29495 32456 29504
rect 32404 29461 32413 29495
rect 32413 29461 32447 29495
rect 32447 29461 32456 29495
rect 32404 29452 32456 29461
rect 33232 29452 33284 29504
rect 4874 29350 4926 29402
rect 4938 29350 4990 29402
rect 5002 29350 5054 29402
rect 5066 29350 5118 29402
rect 5130 29350 5182 29402
rect 35594 29350 35646 29402
rect 35658 29350 35710 29402
rect 35722 29350 35774 29402
rect 35786 29350 35838 29402
rect 35850 29350 35902 29402
rect 9312 29248 9364 29300
rect 6092 29180 6144 29232
rect 7288 29180 7340 29232
rect 8116 29180 8168 29232
rect 11244 29248 11296 29300
rect 14648 29248 14700 29300
rect 13636 29180 13688 29232
rect 15568 29180 15620 29232
rect 6460 29112 6512 29164
rect 11704 29112 11756 29164
rect 9312 29087 9364 29096
rect 9312 29053 9321 29087
rect 9321 29053 9355 29087
rect 9355 29053 9364 29087
rect 9312 29044 9364 29053
rect 11152 29044 11204 29096
rect 12624 29087 12676 29096
rect 11796 29019 11848 29028
rect 11796 28985 11805 29019
rect 11805 28985 11839 29019
rect 11839 28985 11848 29019
rect 11796 28976 11848 28985
rect 12624 29053 12633 29087
rect 12633 29053 12667 29087
rect 12667 29053 12676 29087
rect 12624 29044 12676 29053
rect 14556 29087 14608 29096
rect 14556 29053 14565 29087
rect 14565 29053 14599 29087
rect 14599 29053 14608 29087
rect 14556 29044 14608 29053
rect 15292 29044 15344 29096
rect 18420 29248 18472 29300
rect 21640 29248 21692 29300
rect 23756 29248 23808 29300
rect 26700 29248 26752 29300
rect 29184 29248 29236 29300
rect 29552 29291 29604 29300
rect 29552 29257 29561 29291
rect 29561 29257 29595 29291
rect 29595 29257 29604 29291
rect 29552 29248 29604 29257
rect 29644 29248 29696 29300
rect 31300 29291 31352 29300
rect 31300 29257 31309 29291
rect 31309 29257 31343 29291
rect 31343 29257 31352 29291
rect 31300 29248 31352 29257
rect 31668 29248 31720 29300
rect 32220 29248 32272 29300
rect 33140 29248 33192 29300
rect 26516 29180 26568 29232
rect 30012 29180 30064 29232
rect 19616 29155 19668 29164
rect 19616 29121 19625 29155
rect 19625 29121 19659 29155
rect 19659 29121 19668 29155
rect 19616 29112 19668 29121
rect 20260 29155 20312 29164
rect 20260 29121 20269 29155
rect 20269 29121 20303 29155
rect 20303 29121 20312 29155
rect 20260 29112 20312 29121
rect 22192 29112 22244 29164
rect 23572 29112 23624 29164
rect 27436 29155 27488 29164
rect 27436 29121 27445 29155
rect 27445 29121 27479 29155
rect 27479 29121 27488 29155
rect 27436 29112 27488 29121
rect 28356 29155 28408 29164
rect 28356 29121 28365 29155
rect 28365 29121 28399 29155
rect 28399 29121 28408 29155
rect 28356 29112 28408 29121
rect 28540 29155 28592 29164
rect 28540 29121 28549 29155
rect 28549 29121 28583 29155
rect 28583 29121 28592 29155
rect 28540 29112 28592 29121
rect 28908 29155 28960 29164
rect 28908 29121 28917 29155
rect 28917 29121 28951 29155
rect 28951 29121 28960 29155
rect 28908 29112 28960 29121
rect 18604 29044 18656 29096
rect 18972 29087 19024 29096
rect 18972 29053 18981 29087
rect 18981 29053 19015 29087
rect 19015 29053 19024 29087
rect 18972 29044 19024 29053
rect 21272 29044 21324 29096
rect 22836 29087 22888 29096
rect 22836 29053 22845 29087
rect 22845 29053 22879 29087
rect 22879 29053 22888 29087
rect 22836 29044 22888 29053
rect 8392 28908 8444 28960
rect 9588 28908 9640 28960
rect 13820 28976 13872 29028
rect 14096 28951 14148 28960
rect 14096 28917 14105 28951
rect 14105 28917 14139 28951
rect 14139 28917 14148 28951
rect 14096 28908 14148 28917
rect 16304 28951 16356 28960
rect 16304 28917 16313 28951
rect 16313 28917 16347 28951
rect 16347 28917 16356 28951
rect 16304 28908 16356 28917
rect 22652 28976 22704 29028
rect 23572 28976 23624 29028
rect 24124 29087 24176 29096
rect 24124 29053 24133 29087
rect 24133 29053 24167 29087
rect 24167 29053 24176 29087
rect 24860 29087 24912 29096
rect 24124 29044 24176 29053
rect 24860 29053 24869 29087
rect 24869 29053 24903 29087
rect 24903 29053 24912 29087
rect 24860 29044 24912 29053
rect 25136 29087 25188 29096
rect 25136 29053 25145 29087
rect 25145 29053 25179 29087
rect 25179 29053 25188 29087
rect 25136 29044 25188 29053
rect 28448 29044 28500 29096
rect 28632 29087 28684 29096
rect 28632 29053 28641 29087
rect 28641 29053 28675 29087
rect 28675 29053 28684 29087
rect 28632 29044 28684 29053
rect 22100 28908 22152 28960
rect 26884 28976 26936 29028
rect 28816 29044 28868 29096
rect 29828 29112 29880 29164
rect 32036 29180 32088 29232
rect 31760 29112 31812 29164
rect 34520 29112 34572 29164
rect 30380 29044 30432 29096
rect 33232 29044 33284 29096
rect 34428 29087 34480 29096
rect 34428 29053 34437 29087
rect 34437 29053 34471 29087
rect 34471 29053 34480 29087
rect 34428 29044 34480 29053
rect 29460 28908 29512 28960
rect 32496 28951 32548 28960
rect 32496 28917 32505 28951
rect 32505 28917 32539 28951
rect 32539 28917 32548 28951
rect 32496 28908 32548 28917
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 12624 28704 12676 28756
rect 15568 28747 15620 28756
rect 15568 28713 15577 28747
rect 15577 28713 15611 28747
rect 15611 28713 15620 28747
rect 15568 28704 15620 28713
rect 16120 28704 16172 28756
rect 25136 28704 25188 28756
rect 26516 28747 26568 28756
rect 26516 28713 26525 28747
rect 26525 28713 26559 28747
rect 26559 28713 26568 28747
rect 26516 28704 26568 28713
rect 29000 28747 29052 28756
rect 29000 28713 29009 28747
rect 29009 28713 29043 28747
rect 29043 28713 29052 28747
rect 29000 28704 29052 28713
rect 29092 28704 29144 28756
rect 31300 28704 31352 28756
rect 34520 28704 34572 28756
rect 9496 28636 9548 28688
rect 8208 28568 8260 28620
rect 9588 28611 9640 28620
rect 6828 28364 6880 28416
rect 9588 28577 9597 28611
rect 9597 28577 9631 28611
rect 9631 28577 9640 28611
rect 9588 28568 9640 28577
rect 12532 28568 12584 28620
rect 18144 28636 18196 28688
rect 18236 28568 18288 28620
rect 18420 28568 18472 28620
rect 18696 28611 18748 28620
rect 18696 28577 18705 28611
rect 18705 28577 18739 28611
rect 18739 28577 18748 28611
rect 18696 28568 18748 28577
rect 18972 28568 19024 28620
rect 14188 28500 14240 28552
rect 14648 28500 14700 28552
rect 15476 28543 15528 28552
rect 15476 28509 15485 28543
rect 15485 28509 15519 28543
rect 15519 28509 15528 28543
rect 15476 28500 15528 28509
rect 16856 28500 16908 28552
rect 19892 28500 19944 28552
rect 24124 28568 24176 28620
rect 24952 28568 25004 28620
rect 25136 28568 25188 28620
rect 8300 28364 8352 28416
rect 14832 28432 14884 28484
rect 22836 28500 22888 28552
rect 26884 28636 26936 28688
rect 28356 28568 28408 28620
rect 28724 28568 28776 28620
rect 29184 28636 29236 28688
rect 26608 28543 26660 28552
rect 26608 28509 26617 28543
rect 26617 28509 26651 28543
rect 26651 28509 26660 28543
rect 26608 28500 26660 28509
rect 28264 28543 28316 28552
rect 28264 28509 28273 28543
rect 28273 28509 28307 28543
rect 28307 28509 28316 28543
rect 28264 28500 28316 28509
rect 29644 28568 29696 28620
rect 20812 28432 20864 28484
rect 23480 28432 23532 28484
rect 26884 28432 26936 28484
rect 28908 28500 28960 28552
rect 29828 28543 29880 28552
rect 29828 28509 29837 28543
rect 29837 28509 29871 28543
rect 29871 28509 29880 28543
rect 33232 28611 33284 28620
rect 33232 28577 33241 28611
rect 33241 28577 33275 28611
rect 33275 28577 33284 28611
rect 33232 28568 33284 28577
rect 29828 28500 29880 28509
rect 28540 28432 28592 28484
rect 29276 28432 29328 28484
rect 29460 28432 29512 28484
rect 31944 28500 31996 28552
rect 33140 28500 33192 28552
rect 35072 28543 35124 28552
rect 32404 28432 32456 28484
rect 35072 28509 35081 28543
rect 35081 28509 35115 28543
rect 35115 28509 35124 28543
rect 35072 28500 35124 28509
rect 35440 28500 35492 28552
rect 9220 28364 9272 28416
rect 11244 28407 11296 28416
rect 11244 28373 11253 28407
rect 11253 28373 11287 28407
rect 11287 28373 11296 28407
rect 11244 28364 11296 28373
rect 11336 28407 11388 28416
rect 11336 28373 11345 28407
rect 11345 28373 11379 28407
rect 11379 28373 11388 28407
rect 11336 28364 11388 28373
rect 11888 28364 11940 28416
rect 13544 28407 13596 28416
rect 13544 28373 13553 28407
rect 13553 28373 13587 28407
rect 13587 28373 13596 28407
rect 13544 28364 13596 28373
rect 14648 28407 14700 28416
rect 14648 28373 14657 28407
rect 14657 28373 14691 28407
rect 14691 28373 14700 28407
rect 14648 28364 14700 28373
rect 14740 28407 14792 28416
rect 14740 28373 14749 28407
rect 14749 28373 14783 28407
rect 14783 28373 14792 28407
rect 16120 28407 16172 28416
rect 14740 28364 14792 28373
rect 16120 28373 16129 28407
rect 16129 28373 16163 28407
rect 16163 28373 16172 28407
rect 16120 28364 16172 28373
rect 17592 28364 17644 28416
rect 18052 28364 18104 28416
rect 18420 28364 18472 28416
rect 19984 28364 20036 28416
rect 20536 28364 20588 28416
rect 23204 28407 23256 28416
rect 23204 28373 23213 28407
rect 23213 28373 23247 28407
rect 23247 28373 23256 28407
rect 23204 28364 23256 28373
rect 24584 28364 24636 28416
rect 29920 28364 29972 28416
rect 31024 28364 31076 28416
rect 31208 28364 31260 28416
rect 33416 28364 33468 28416
rect 34612 28364 34664 28416
rect 35164 28364 35216 28416
rect 4874 28262 4926 28314
rect 4938 28262 4990 28314
rect 5002 28262 5054 28314
rect 5066 28262 5118 28314
rect 5130 28262 5182 28314
rect 35594 28262 35646 28314
rect 35658 28262 35710 28314
rect 35722 28262 35774 28314
rect 35786 28262 35838 28314
rect 35850 28262 35902 28314
rect 1860 28024 1912 28076
rect 7104 28160 7156 28212
rect 8300 28203 8352 28212
rect 6828 28135 6880 28144
rect 6828 28101 6837 28135
rect 6837 28101 6871 28135
rect 6871 28101 6880 28135
rect 6828 28092 6880 28101
rect 7288 28092 7340 28144
rect 8300 28169 8309 28203
rect 8309 28169 8343 28203
rect 8343 28169 8352 28203
rect 8300 28160 8352 28169
rect 11244 28160 11296 28212
rect 11336 28160 11388 28212
rect 14188 28203 14240 28212
rect 14188 28169 14197 28203
rect 14197 28169 14231 28203
rect 14231 28169 14240 28203
rect 14188 28160 14240 28169
rect 14648 28160 14700 28212
rect 16856 28203 16908 28212
rect 16856 28169 16865 28203
rect 16865 28169 16899 28203
rect 16899 28169 16908 28203
rect 16856 28160 16908 28169
rect 14096 28092 14148 28144
rect 8760 28067 8812 28076
rect 8760 28033 8769 28067
rect 8769 28033 8803 28067
rect 8803 28033 8812 28067
rect 8760 28024 8812 28033
rect 11888 28067 11940 28076
rect 9312 27956 9364 28008
rect 11888 28033 11897 28067
rect 11897 28033 11931 28067
rect 11931 28033 11940 28067
rect 11888 28024 11940 28033
rect 13084 28024 13136 28076
rect 13728 28024 13780 28076
rect 14740 28092 14792 28144
rect 16304 28092 16356 28144
rect 12716 27956 12768 28008
rect 17592 28024 17644 28076
rect 18052 28067 18104 28076
rect 18052 28033 18061 28067
rect 18061 28033 18095 28067
rect 18095 28033 18104 28067
rect 18052 28024 18104 28033
rect 18696 28092 18748 28144
rect 20812 28160 20864 28212
rect 28264 28160 28316 28212
rect 29920 28160 29972 28212
rect 19984 28092 20036 28144
rect 22284 28092 22336 28144
rect 24768 28092 24820 28144
rect 22100 28024 22152 28076
rect 22192 28067 22244 28076
rect 22192 28033 22201 28067
rect 22201 28033 22235 28067
rect 22235 28033 22244 28067
rect 23020 28067 23072 28076
rect 22192 28024 22244 28033
rect 23020 28033 23029 28067
rect 23029 28033 23063 28067
rect 23063 28033 23072 28067
rect 23020 28024 23072 28033
rect 24216 28067 24268 28076
rect 24216 28033 24225 28067
rect 24225 28033 24259 28067
rect 24259 28033 24268 28067
rect 24216 28024 24268 28033
rect 15016 27888 15068 27940
rect 18236 27888 18288 27940
rect 1584 27863 1636 27872
rect 1584 27829 1593 27863
rect 1593 27829 1627 27863
rect 1627 27829 1636 27863
rect 1584 27820 1636 27829
rect 13636 27863 13688 27872
rect 13636 27829 13645 27863
rect 13645 27829 13679 27863
rect 13679 27829 13688 27863
rect 13636 27820 13688 27829
rect 24124 27956 24176 28008
rect 25136 27999 25188 28008
rect 25136 27965 25145 27999
rect 25145 27965 25179 27999
rect 25179 27965 25188 27999
rect 25136 27956 25188 27965
rect 26608 28024 26660 28076
rect 28816 28024 28868 28076
rect 30748 28160 30800 28212
rect 33508 28160 33560 28212
rect 32496 28092 32548 28144
rect 32956 28092 33008 28144
rect 28908 27956 28960 28008
rect 31116 28024 31168 28076
rect 31576 28024 31628 28076
rect 35072 28160 35124 28212
rect 30564 27956 30616 28008
rect 31392 27956 31444 28008
rect 31944 27956 31996 28008
rect 34428 28092 34480 28144
rect 35164 28135 35216 28144
rect 30472 27888 30524 27940
rect 33324 27888 33376 27940
rect 18972 27820 19024 27872
rect 19708 27820 19760 27872
rect 20444 27863 20496 27872
rect 20444 27829 20453 27863
rect 20453 27829 20487 27863
rect 20487 27829 20496 27863
rect 20444 27820 20496 27829
rect 22100 27863 22152 27872
rect 22100 27829 22109 27863
rect 22109 27829 22143 27863
rect 22143 27829 22152 27863
rect 23848 27863 23900 27872
rect 22100 27820 22152 27829
rect 23848 27829 23857 27863
rect 23857 27829 23891 27863
rect 23891 27829 23900 27863
rect 23848 27820 23900 27829
rect 26148 27820 26200 27872
rect 27528 27820 27580 27872
rect 29184 27863 29236 27872
rect 29184 27829 29193 27863
rect 29193 27829 29227 27863
rect 29227 27829 29236 27863
rect 29184 27820 29236 27829
rect 29828 27820 29880 27872
rect 32036 27820 32088 27872
rect 35164 28101 35173 28135
rect 35173 28101 35207 28135
rect 35207 28101 35216 28135
rect 35164 28092 35216 28101
rect 36176 28092 36228 28144
rect 36636 27863 36688 27872
rect 36636 27829 36645 27863
rect 36645 27829 36679 27863
rect 36679 27829 36688 27863
rect 36636 27820 36688 27829
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 16120 27659 16172 27668
rect 16120 27625 16150 27659
rect 16150 27625 16172 27659
rect 16120 27616 16172 27625
rect 22192 27616 22244 27668
rect 7288 27591 7340 27600
rect 7288 27557 7297 27591
rect 7297 27557 7331 27591
rect 7331 27557 7340 27591
rect 7288 27548 7340 27557
rect 14556 27548 14608 27600
rect 8208 27480 8260 27532
rect 9312 27480 9364 27532
rect 11060 27480 11112 27532
rect 12164 27480 12216 27532
rect 12348 27480 12400 27532
rect 12532 27480 12584 27532
rect 18512 27548 18564 27600
rect 18236 27523 18288 27532
rect 18236 27489 18245 27523
rect 18245 27489 18279 27523
rect 18279 27489 18288 27523
rect 18236 27480 18288 27489
rect 18420 27523 18472 27532
rect 18420 27489 18429 27523
rect 18429 27489 18463 27523
rect 18463 27489 18472 27523
rect 20444 27548 20496 27600
rect 18420 27480 18472 27489
rect 20812 27548 20864 27600
rect 23480 27591 23532 27600
rect 23480 27557 23489 27591
rect 23489 27557 23523 27591
rect 23523 27557 23532 27591
rect 23480 27548 23532 27557
rect 8760 27412 8812 27464
rect 9588 27455 9640 27464
rect 9588 27421 9597 27455
rect 9597 27421 9631 27455
rect 9631 27421 9640 27455
rect 9588 27412 9640 27421
rect 14556 27455 14608 27464
rect 14556 27421 14565 27455
rect 14565 27421 14599 27455
rect 14599 27421 14608 27455
rect 14556 27412 14608 27421
rect 9680 27344 9732 27396
rect 7932 27276 7984 27328
rect 9220 27276 9272 27328
rect 11796 27344 11848 27396
rect 12348 27344 12400 27396
rect 13728 27344 13780 27396
rect 19340 27412 19392 27464
rect 21272 27455 21324 27464
rect 11152 27276 11204 27328
rect 13084 27319 13136 27328
rect 13084 27285 13093 27319
rect 13093 27285 13127 27319
rect 13127 27285 13136 27319
rect 13084 27276 13136 27285
rect 14188 27276 14240 27328
rect 18880 27344 18932 27396
rect 21272 27421 21281 27455
rect 21281 27421 21315 27455
rect 21315 27421 21324 27455
rect 21272 27412 21324 27421
rect 23204 27412 23256 27464
rect 23480 27412 23532 27464
rect 28816 27616 28868 27668
rect 35440 27616 35492 27668
rect 31760 27548 31812 27600
rect 23664 27480 23716 27532
rect 24860 27480 24912 27532
rect 34612 27548 34664 27600
rect 36176 27591 36228 27600
rect 36176 27557 36185 27591
rect 36185 27557 36219 27591
rect 36219 27557 36228 27591
rect 36176 27548 36228 27557
rect 37096 27591 37148 27600
rect 37096 27557 37105 27591
rect 37105 27557 37139 27591
rect 37139 27557 37148 27591
rect 37096 27548 37148 27557
rect 32496 27523 32548 27532
rect 32496 27489 32505 27523
rect 32505 27489 32539 27523
rect 32539 27489 32548 27523
rect 32496 27480 32548 27489
rect 33324 27480 33376 27532
rect 24676 27412 24728 27464
rect 27160 27455 27212 27464
rect 27160 27421 27169 27455
rect 27169 27421 27203 27455
rect 27203 27421 27212 27455
rect 27160 27412 27212 27421
rect 24952 27344 25004 27396
rect 25228 27387 25280 27396
rect 25228 27353 25237 27387
rect 25237 27353 25271 27387
rect 25271 27353 25280 27387
rect 25228 27344 25280 27353
rect 26884 27344 26936 27396
rect 27436 27387 27488 27396
rect 27436 27353 27445 27387
rect 27445 27353 27479 27387
rect 27479 27353 27488 27387
rect 27436 27344 27488 27353
rect 27528 27344 27580 27396
rect 31024 27412 31076 27464
rect 31392 27455 31444 27464
rect 31392 27421 31401 27455
rect 31401 27421 31435 27455
rect 31435 27421 31444 27455
rect 31392 27412 31444 27421
rect 31576 27344 31628 27396
rect 16488 27276 16540 27328
rect 17592 27319 17644 27328
rect 17592 27285 17601 27319
rect 17601 27285 17635 27319
rect 17635 27285 17644 27319
rect 17592 27276 17644 27285
rect 18420 27276 18472 27328
rect 19432 27319 19484 27328
rect 19432 27285 19441 27319
rect 19441 27285 19475 27319
rect 19475 27285 19484 27319
rect 19432 27276 19484 27285
rect 20628 27319 20680 27328
rect 20628 27285 20637 27319
rect 20637 27285 20671 27319
rect 20671 27285 20680 27319
rect 20628 27276 20680 27285
rect 21364 27319 21416 27328
rect 21364 27285 21373 27319
rect 21373 27285 21407 27319
rect 21407 27285 21416 27319
rect 21364 27276 21416 27285
rect 22192 27319 22244 27328
rect 22192 27285 22201 27319
rect 22201 27285 22235 27319
rect 22235 27285 22244 27319
rect 22192 27276 22244 27285
rect 22652 27319 22704 27328
rect 22652 27285 22661 27319
rect 22661 27285 22695 27319
rect 22695 27285 22704 27319
rect 22652 27276 22704 27285
rect 24584 27276 24636 27328
rect 28356 27276 28408 27328
rect 30748 27319 30800 27328
rect 30748 27285 30757 27319
rect 30757 27285 30791 27319
rect 30791 27285 30800 27319
rect 30748 27276 30800 27285
rect 30840 27276 30892 27328
rect 32864 27412 32916 27464
rect 34796 27480 34848 27532
rect 35164 27480 35216 27532
rect 36636 27480 36688 27532
rect 33048 27344 33100 27396
rect 36360 27412 36412 27464
rect 37004 27412 37056 27464
rect 32864 27276 32916 27328
rect 35164 27319 35216 27328
rect 35164 27285 35173 27319
rect 35173 27285 35207 27319
rect 35207 27285 35216 27319
rect 35164 27276 35216 27285
rect 36452 27276 36504 27328
rect 4874 27174 4926 27226
rect 4938 27174 4990 27226
rect 5002 27174 5054 27226
rect 5066 27174 5118 27226
rect 5130 27174 5182 27226
rect 35594 27174 35646 27226
rect 35658 27174 35710 27226
rect 35722 27174 35774 27226
rect 35786 27174 35838 27226
rect 35850 27174 35902 27226
rect 9220 27072 9272 27124
rect 9588 27115 9640 27124
rect 9588 27081 9597 27115
rect 9597 27081 9631 27115
rect 9631 27081 9640 27115
rect 9588 27072 9640 27081
rect 9680 27072 9732 27124
rect 12164 27115 12216 27124
rect 12164 27081 12173 27115
rect 12173 27081 12207 27115
rect 12207 27081 12216 27115
rect 12164 27072 12216 27081
rect 8392 27004 8444 27056
rect 11244 27004 11296 27056
rect 12348 27004 12400 27056
rect 11060 26936 11112 26988
rect 11704 26936 11756 26988
rect 13728 27072 13780 27124
rect 14556 27072 14608 27124
rect 13544 27047 13596 27056
rect 13544 27013 13553 27047
rect 13553 27013 13587 27047
rect 13587 27013 13596 27047
rect 13544 27004 13596 27013
rect 13636 27004 13688 27056
rect 16764 27004 16816 27056
rect 21364 27072 21416 27124
rect 22652 27072 22704 27124
rect 24216 27072 24268 27124
rect 20628 27004 20680 27056
rect 7748 26868 7800 26920
rect 9036 26732 9088 26784
rect 11428 26732 11480 26784
rect 12716 26868 12768 26920
rect 15016 26911 15068 26920
rect 11796 26800 11848 26852
rect 15016 26877 15025 26911
rect 15025 26877 15059 26911
rect 15059 26877 15068 26911
rect 15016 26868 15068 26877
rect 20076 26936 20128 26988
rect 20720 26936 20772 26988
rect 23664 27047 23716 27056
rect 23664 27013 23673 27047
rect 23673 27013 23707 27047
rect 23707 27013 23716 27047
rect 23664 27004 23716 27013
rect 24584 27004 24636 27056
rect 22192 26979 22244 26988
rect 22192 26945 22201 26979
rect 22201 26945 22235 26979
rect 22235 26945 22244 26979
rect 25228 27072 25280 27124
rect 27436 27072 27488 27124
rect 29184 27072 29236 27124
rect 30748 27115 30800 27124
rect 30748 27081 30757 27115
rect 30757 27081 30791 27115
rect 30791 27081 30800 27115
rect 30748 27072 30800 27081
rect 28632 27004 28684 27056
rect 32956 27072 33008 27124
rect 33324 27072 33376 27124
rect 22192 26936 22244 26945
rect 26148 26936 26200 26988
rect 26700 26936 26752 26988
rect 28356 26979 28408 26988
rect 28356 26945 28365 26979
rect 28365 26945 28399 26979
rect 28399 26945 28408 26979
rect 28356 26936 28408 26945
rect 28540 26979 28592 26988
rect 28540 26945 28549 26979
rect 28549 26945 28583 26979
rect 28583 26945 28592 26979
rect 28540 26936 28592 26945
rect 15108 26800 15160 26852
rect 18972 26868 19024 26920
rect 19708 26911 19760 26920
rect 19708 26877 19717 26911
rect 19717 26877 19751 26911
rect 19751 26877 19760 26911
rect 19708 26868 19760 26877
rect 17408 26800 17460 26852
rect 19800 26800 19852 26852
rect 25136 26868 25188 26920
rect 26608 26868 26660 26920
rect 27344 26911 27396 26920
rect 27344 26877 27353 26911
rect 27353 26877 27387 26911
rect 27387 26877 27396 26911
rect 30472 26936 30524 26988
rect 31392 27004 31444 27056
rect 30564 26911 30616 26920
rect 27344 26868 27396 26877
rect 30564 26877 30573 26911
rect 30573 26877 30607 26911
rect 30607 26877 30616 26911
rect 30564 26868 30616 26877
rect 28540 26800 28592 26852
rect 30840 26800 30892 26852
rect 32312 26936 32364 26988
rect 33508 27004 33560 27056
rect 32956 26868 33008 26920
rect 34244 26936 34296 26988
rect 35808 26979 35860 26988
rect 35808 26945 35817 26979
rect 35817 26945 35851 26979
rect 35851 26945 35860 26979
rect 35808 26936 35860 26945
rect 36452 26979 36504 26988
rect 36452 26945 36461 26979
rect 36461 26945 36495 26979
rect 36495 26945 36504 26979
rect 36452 26936 36504 26945
rect 32496 26800 32548 26852
rect 12532 26732 12584 26784
rect 17224 26732 17276 26784
rect 18420 26732 18472 26784
rect 19616 26732 19668 26784
rect 19892 26732 19944 26784
rect 20996 26732 21048 26784
rect 22376 26732 22428 26784
rect 28448 26732 28500 26784
rect 29276 26775 29328 26784
rect 29276 26741 29285 26775
rect 29285 26741 29319 26775
rect 29319 26741 29328 26775
rect 29276 26732 29328 26741
rect 31668 26732 31720 26784
rect 32956 26732 33008 26784
rect 33968 26732 34020 26784
rect 34796 26868 34848 26920
rect 34612 26800 34664 26852
rect 34704 26800 34756 26852
rect 34796 26732 34848 26784
rect 35440 26732 35492 26784
rect 35624 26732 35676 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 7748 26571 7800 26580
rect 7748 26537 7757 26571
rect 7757 26537 7791 26571
rect 7791 26537 7800 26571
rect 7748 26528 7800 26537
rect 8392 26528 8444 26580
rect 18328 26528 18380 26580
rect 18880 26571 18932 26580
rect 18880 26537 18889 26571
rect 18889 26537 18923 26571
rect 18923 26537 18932 26571
rect 18880 26528 18932 26537
rect 18972 26528 19024 26580
rect 22376 26528 22428 26580
rect 22652 26528 22704 26580
rect 24952 26528 25004 26580
rect 10048 26460 10100 26512
rect 10508 26460 10560 26512
rect 7932 26367 7984 26376
rect 7932 26333 7941 26367
rect 7941 26333 7975 26367
rect 7975 26333 7984 26367
rect 7932 26324 7984 26333
rect 8760 26324 8812 26376
rect 10048 26367 10100 26376
rect 10048 26333 10057 26367
rect 10057 26333 10091 26367
rect 10091 26333 10100 26367
rect 10048 26324 10100 26333
rect 11244 26392 11296 26444
rect 11796 26435 11848 26444
rect 11796 26401 11805 26435
rect 11805 26401 11839 26435
rect 11839 26401 11848 26435
rect 11796 26392 11848 26401
rect 13084 26392 13136 26444
rect 15108 26435 15160 26444
rect 15108 26401 15117 26435
rect 15117 26401 15151 26435
rect 15151 26401 15160 26435
rect 15108 26392 15160 26401
rect 11152 26367 11204 26376
rect 11152 26333 11161 26367
rect 11161 26333 11195 26367
rect 11195 26333 11204 26367
rect 11152 26324 11204 26333
rect 19800 26460 19852 26512
rect 19892 26460 19944 26512
rect 17408 26435 17460 26444
rect 17408 26401 17417 26435
rect 17417 26401 17451 26435
rect 17451 26401 17460 26435
rect 17408 26392 17460 26401
rect 17592 26324 17644 26376
rect 18236 26435 18288 26444
rect 18236 26401 18245 26435
rect 18245 26401 18279 26435
rect 18279 26401 18288 26435
rect 18236 26392 18288 26401
rect 18420 26435 18472 26444
rect 18420 26401 18429 26435
rect 18429 26401 18463 26435
rect 18463 26401 18472 26435
rect 18420 26392 18472 26401
rect 20628 26392 20680 26444
rect 23664 26460 23716 26512
rect 26884 26528 26936 26580
rect 28448 26528 28500 26580
rect 30472 26528 30524 26580
rect 32312 26528 32364 26580
rect 34244 26571 34296 26580
rect 34244 26537 34253 26571
rect 34253 26537 34287 26571
rect 34287 26537 34296 26571
rect 34244 26528 34296 26537
rect 35808 26528 35860 26580
rect 23480 26392 23532 26444
rect 23756 26392 23808 26444
rect 22100 26324 22152 26376
rect 23848 26324 23900 26376
rect 24676 26392 24728 26444
rect 26240 26392 26292 26444
rect 30656 26460 30708 26512
rect 31668 26435 31720 26444
rect 27344 26324 27396 26376
rect 31668 26401 31677 26435
rect 31677 26401 31711 26435
rect 31711 26401 31720 26435
rect 31668 26392 31720 26401
rect 33416 26460 33468 26512
rect 11336 26256 11388 26308
rect 11428 26256 11480 26308
rect 20996 26299 21048 26308
rect 9680 26231 9732 26240
rect 9680 26197 9689 26231
rect 9689 26197 9723 26231
rect 9723 26197 9732 26231
rect 9680 26188 9732 26197
rect 10140 26231 10192 26240
rect 10140 26197 10149 26231
rect 10149 26197 10183 26231
rect 10183 26197 10192 26231
rect 10140 26188 10192 26197
rect 13820 26188 13872 26240
rect 18512 26231 18564 26240
rect 18512 26197 18521 26231
rect 18521 26197 18555 26231
rect 18555 26197 18564 26231
rect 19524 26231 19576 26240
rect 18512 26188 18564 26197
rect 19524 26197 19533 26231
rect 19533 26197 19567 26231
rect 19567 26197 19576 26231
rect 19524 26188 19576 26197
rect 19892 26231 19944 26240
rect 19892 26197 19901 26231
rect 19901 26197 19935 26231
rect 19935 26197 19944 26231
rect 19892 26188 19944 26197
rect 20996 26265 21005 26299
rect 21005 26265 21039 26299
rect 21039 26265 21048 26299
rect 20996 26256 21048 26265
rect 25320 26299 25372 26308
rect 23480 26231 23532 26240
rect 23480 26197 23489 26231
rect 23489 26197 23523 26231
rect 23523 26197 23532 26231
rect 23480 26188 23532 26197
rect 24584 26231 24636 26240
rect 24584 26197 24593 26231
rect 24593 26197 24627 26231
rect 24627 26197 24636 26231
rect 24584 26188 24636 26197
rect 25320 26265 25329 26299
rect 25329 26265 25363 26299
rect 25363 26265 25372 26299
rect 25320 26256 25372 26265
rect 28632 26324 28684 26376
rect 31944 26367 31996 26376
rect 31944 26333 31953 26367
rect 31953 26333 31987 26367
rect 31987 26333 31996 26367
rect 33048 26392 33100 26444
rect 33876 26435 33928 26444
rect 33876 26401 33885 26435
rect 33885 26401 33919 26435
rect 33919 26401 33928 26435
rect 33876 26392 33928 26401
rect 32956 26367 33008 26376
rect 31944 26324 31996 26333
rect 28540 26299 28592 26308
rect 28540 26265 28549 26299
rect 28549 26265 28583 26299
rect 28583 26265 28592 26299
rect 28540 26256 28592 26265
rect 31208 26256 31260 26308
rect 32956 26333 32965 26367
rect 32965 26333 32999 26367
rect 32999 26333 33008 26367
rect 32956 26324 33008 26333
rect 26056 26188 26108 26240
rect 26332 26188 26384 26240
rect 27712 26231 27764 26240
rect 27712 26197 27721 26231
rect 27721 26197 27755 26231
rect 27755 26197 27764 26231
rect 27712 26188 27764 26197
rect 28908 26231 28960 26240
rect 28908 26197 28917 26231
rect 28917 26197 28951 26231
rect 28951 26197 28960 26231
rect 28908 26188 28960 26197
rect 31300 26188 31352 26240
rect 32588 26256 32640 26308
rect 33140 26367 33192 26376
rect 33140 26333 33149 26367
rect 33149 26333 33183 26367
rect 33183 26333 33192 26367
rect 33968 26367 34020 26376
rect 33140 26324 33192 26333
rect 33968 26333 33977 26367
rect 33977 26333 34011 26367
rect 34011 26333 34020 26367
rect 33968 26324 34020 26333
rect 34612 26460 34664 26512
rect 34520 26392 34572 26444
rect 35624 26435 35676 26444
rect 35624 26401 35633 26435
rect 35633 26401 35667 26435
rect 35667 26401 35676 26435
rect 35624 26392 35676 26401
rect 35348 26324 35400 26376
rect 34520 26256 34572 26308
rect 36452 26256 36504 26308
rect 33692 26188 33744 26240
rect 4874 26086 4926 26138
rect 4938 26086 4990 26138
rect 5002 26086 5054 26138
rect 5066 26086 5118 26138
rect 5130 26086 5182 26138
rect 35594 26086 35646 26138
rect 35658 26086 35710 26138
rect 35722 26086 35774 26138
rect 35786 26086 35838 26138
rect 35850 26086 35902 26138
rect 9128 25848 9180 25900
rect 9772 25916 9824 25968
rect 9956 25916 10008 25968
rect 12808 25984 12860 26036
rect 14188 25959 14240 25968
rect 14188 25925 14197 25959
rect 14197 25925 14231 25959
rect 14231 25925 14240 25959
rect 14188 25916 14240 25925
rect 15200 25916 15252 25968
rect 18328 25959 18380 25968
rect 18328 25925 18337 25959
rect 18337 25925 18371 25959
rect 18371 25925 18380 25959
rect 18328 25916 18380 25925
rect 19708 25984 19760 26036
rect 20996 25916 21048 25968
rect 10876 25848 10928 25900
rect 13820 25848 13872 25900
rect 8576 25780 8628 25832
rect 13728 25780 13780 25832
rect 10508 25712 10560 25764
rect 15660 25780 15712 25832
rect 17224 25848 17276 25900
rect 19524 25848 19576 25900
rect 23756 25984 23808 26036
rect 26056 26027 26108 26036
rect 26056 25993 26065 26027
rect 26065 25993 26099 26027
rect 26099 25993 26108 26027
rect 26056 25984 26108 25993
rect 28356 25984 28408 26036
rect 25320 25916 25372 25968
rect 24768 25848 24820 25900
rect 26332 25916 26384 25968
rect 27712 25916 27764 25968
rect 27896 25916 27948 25968
rect 32036 25984 32088 26036
rect 33876 25984 33928 26036
rect 18604 25823 18656 25832
rect 18604 25789 18613 25823
rect 18613 25789 18647 25823
rect 18647 25789 18656 25823
rect 19708 25823 19760 25832
rect 18604 25780 18656 25789
rect 19708 25789 19717 25823
rect 19717 25789 19751 25823
rect 19751 25789 19760 25823
rect 19708 25780 19760 25789
rect 24584 25780 24636 25832
rect 19432 25712 19484 25764
rect 23480 25712 23532 25764
rect 25596 25780 25648 25832
rect 8484 25687 8536 25696
rect 8484 25653 8493 25687
rect 8493 25653 8527 25687
rect 8527 25653 8536 25687
rect 8484 25644 8536 25653
rect 12164 25644 12216 25696
rect 14556 25644 14608 25696
rect 16304 25687 16356 25696
rect 16304 25653 16313 25687
rect 16313 25653 16347 25687
rect 16347 25653 16356 25687
rect 16304 25644 16356 25653
rect 16580 25644 16632 25696
rect 19984 25644 20036 25696
rect 21088 25644 21140 25696
rect 24492 25687 24544 25696
rect 24492 25653 24501 25687
rect 24501 25653 24535 25687
rect 24535 25653 24544 25687
rect 24492 25644 24544 25653
rect 24952 25644 25004 25696
rect 27160 25823 27212 25832
rect 27160 25789 27169 25823
rect 27169 25789 27203 25823
rect 27203 25789 27212 25823
rect 27160 25780 27212 25789
rect 29736 25848 29788 25900
rect 30472 25848 30524 25900
rect 31576 25916 31628 25968
rect 30656 25891 30708 25900
rect 30656 25857 30665 25891
rect 30665 25857 30699 25891
rect 30699 25857 30708 25891
rect 31116 25891 31168 25900
rect 30656 25848 30708 25857
rect 31116 25857 31125 25891
rect 31125 25857 31159 25891
rect 31159 25857 31168 25891
rect 31116 25848 31168 25857
rect 31300 25891 31352 25900
rect 31300 25857 31309 25891
rect 31309 25857 31343 25891
rect 31343 25857 31352 25891
rect 31300 25848 31352 25857
rect 33048 25916 33100 25968
rect 36268 25916 36320 25968
rect 32588 25891 32640 25900
rect 32588 25857 32597 25891
rect 32597 25857 32631 25891
rect 32631 25857 32640 25891
rect 32588 25848 32640 25857
rect 31760 25780 31812 25832
rect 33140 25848 33192 25900
rect 33324 25891 33376 25900
rect 33324 25857 33333 25891
rect 33333 25857 33367 25891
rect 33367 25857 33376 25891
rect 33324 25848 33376 25857
rect 34612 25848 34664 25900
rect 36176 25823 36228 25832
rect 36176 25789 36185 25823
rect 36185 25789 36219 25823
rect 36219 25789 36228 25823
rect 36176 25780 36228 25789
rect 32404 25712 32456 25764
rect 34520 25712 34572 25764
rect 29000 25644 29052 25696
rect 29368 25687 29420 25696
rect 29368 25653 29377 25687
rect 29377 25653 29411 25687
rect 29411 25653 29420 25687
rect 29368 25644 29420 25653
rect 30380 25644 30432 25696
rect 32772 25687 32824 25696
rect 32772 25653 32781 25687
rect 32781 25653 32815 25687
rect 32815 25653 32824 25687
rect 32772 25644 32824 25653
rect 35440 25644 35492 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 8576 25483 8628 25492
rect 8576 25449 8585 25483
rect 8585 25449 8619 25483
rect 8619 25449 8628 25483
rect 8576 25440 8628 25449
rect 12072 25440 12124 25492
rect 18512 25440 18564 25492
rect 20996 25440 21048 25492
rect 28356 25483 28408 25492
rect 28356 25449 28365 25483
rect 28365 25449 28399 25483
rect 28399 25449 28408 25483
rect 28356 25440 28408 25449
rect 29736 25440 29788 25492
rect 31116 25440 31168 25492
rect 31484 25483 31536 25492
rect 31484 25449 31493 25483
rect 31493 25449 31527 25483
rect 31527 25449 31536 25483
rect 31484 25440 31536 25449
rect 31760 25483 31812 25492
rect 31760 25449 31769 25483
rect 31769 25449 31803 25483
rect 31803 25449 31812 25483
rect 31760 25440 31812 25449
rect 32588 25483 32640 25492
rect 32588 25449 32597 25483
rect 32597 25449 32631 25483
rect 32631 25449 32640 25483
rect 32588 25440 32640 25449
rect 36176 25440 36228 25492
rect 36268 25440 36320 25492
rect 19340 25372 19392 25424
rect 9588 25304 9640 25356
rect 11152 25347 11204 25356
rect 11152 25313 11161 25347
rect 11161 25313 11195 25347
rect 11195 25313 11204 25347
rect 11152 25304 11204 25313
rect 14556 25347 14608 25356
rect 14556 25313 14565 25347
rect 14565 25313 14599 25347
rect 14599 25313 14608 25347
rect 14556 25304 14608 25313
rect 14648 25304 14700 25356
rect 7932 25279 7984 25288
rect 7932 25245 7941 25279
rect 7941 25245 7975 25279
rect 7975 25245 7984 25279
rect 7932 25236 7984 25245
rect 9680 25236 9732 25288
rect 10968 25236 11020 25288
rect 13728 25236 13780 25288
rect 16304 25304 16356 25356
rect 19892 25347 19944 25356
rect 19892 25313 19901 25347
rect 19901 25313 19935 25347
rect 19935 25313 19944 25347
rect 19892 25304 19944 25313
rect 20168 25304 20220 25356
rect 23756 25347 23808 25356
rect 23756 25313 23765 25347
rect 23765 25313 23799 25347
rect 23799 25313 23808 25347
rect 23756 25304 23808 25313
rect 23848 25347 23900 25356
rect 23848 25313 23857 25347
rect 23857 25313 23891 25347
rect 23891 25313 23900 25347
rect 23848 25304 23900 25313
rect 26976 25304 27028 25356
rect 30564 25347 30616 25356
rect 30564 25313 30573 25347
rect 30573 25313 30607 25347
rect 30607 25313 30616 25347
rect 30564 25304 30616 25313
rect 30656 25304 30708 25356
rect 8208 25168 8260 25220
rect 7748 25143 7800 25152
rect 7748 25109 7757 25143
rect 7757 25109 7791 25143
rect 7791 25109 7800 25143
rect 7748 25100 7800 25109
rect 9312 25143 9364 25152
rect 9312 25109 9321 25143
rect 9321 25109 9355 25143
rect 9355 25109 9364 25143
rect 9312 25100 9364 25109
rect 10508 25100 10560 25152
rect 12164 25168 12216 25220
rect 14648 25168 14700 25220
rect 15292 25168 15344 25220
rect 17960 25236 18012 25288
rect 20720 25236 20772 25288
rect 16948 25168 17000 25220
rect 14372 25100 14424 25152
rect 15936 25100 15988 25152
rect 19800 25143 19852 25152
rect 19800 25109 19809 25143
rect 19809 25109 19843 25143
rect 19843 25109 19852 25143
rect 19800 25100 19852 25109
rect 22284 25100 22336 25152
rect 24492 25236 24544 25288
rect 24952 25279 25004 25288
rect 24952 25245 24961 25279
rect 24961 25245 24995 25279
rect 24995 25245 25004 25279
rect 24952 25236 25004 25245
rect 24676 25168 24728 25220
rect 29368 25236 29420 25288
rect 29736 25279 29788 25288
rect 29736 25245 29745 25279
rect 29745 25245 29779 25279
rect 29779 25245 29788 25279
rect 29736 25236 29788 25245
rect 30380 25279 30432 25288
rect 30380 25245 30389 25279
rect 30389 25245 30423 25279
rect 30423 25245 30432 25279
rect 30380 25236 30432 25245
rect 31392 25279 31444 25288
rect 26884 25211 26936 25220
rect 26884 25177 26893 25211
rect 26893 25177 26927 25211
rect 26927 25177 26936 25211
rect 26884 25168 26936 25177
rect 29276 25168 29328 25220
rect 31392 25245 31401 25279
rect 31401 25245 31435 25279
rect 31435 25245 31444 25279
rect 31392 25236 31444 25245
rect 33048 25236 33100 25288
rect 34244 25279 34296 25288
rect 34244 25245 34253 25279
rect 34253 25245 34287 25279
rect 34287 25245 34296 25279
rect 34244 25236 34296 25245
rect 32312 25168 32364 25220
rect 33232 25211 33284 25220
rect 33232 25177 33241 25211
rect 33241 25177 33275 25211
rect 33275 25177 33284 25211
rect 33232 25168 33284 25177
rect 33692 25168 33744 25220
rect 34152 25211 34204 25220
rect 34152 25177 34161 25211
rect 34161 25177 34195 25211
rect 34195 25177 34204 25211
rect 35532 25236 35584 25288
rect 36360 25279 36412 25288
rect 36360 25245 36369 25279
rect 36369 25245 36403 25279
rect 36403 25245 36412 25279
rect 36360 25236 36412 25245
rect 34152 25168 34204 25177
rect 24492 25100 24544 25152
rect 24860 25143 24912 25152
rect 24860 25109 24869 25143
rect 24869 25109 24903 25143
rect 24903 25109 24912 25143
rect 24860 25100 24912 25109
rect 25688 25100 25740 25152
rect 25872 25143 25924 25152
rect 25872 25109 25881 25143
rect 25881 25109 25915 25143
rect 25915 25109 25924 25143
rect 25872 25100 25924 25109
rect 30380 25100 30432 25152
rect 34244 25100 34296 25152
rect 34796 25100 34848 25152
rect 4874 24998 4926 25050
rect 4938 24998 4990 25050
rect 5002 24998 5054 25050
rect 5066 24998 5118 25050
rect 5130 24998 5182 25050
rect 35594 24998 35646 25050
rect 35658 24998 35710 25050
rect 35722 24998 35774 25050
rect 35786 24998 35838 25050
rect 35850 24998 35902 25050
rect 10692 24939 10744 24948
rect 10692 24905 10701 24939
rect 10701 24905 10735 24939
rect 10735 24905 10744 24939
rect 12072 24939 12124 24948
rect 10692 24896 10744 24905
rect 12072 24905 12081 24939
rect 12081 24905 12115 24939
rect 12115 24905 12124 24939
rect 12072 24896 12124 24905
rect 21088 24939 21140 24948
rect 21088 24905 21097 24939
rect 21097 24905 21131 24939
rect 21131 24905 21140 24939
rect 21088 24896 21140 24905
rect 23756 24939 23808 24948
rect 23756 24905 23765 24939
rect 23765 24905 23799 24939
rect 23799 24905 23808 24939
rect 23756 24896 23808 24905
rect 24860 24896 24912 24948
rect 25504 24896 25556 24948
rect 26884 24896 26936 24948
rect 28908 24896 28960 24948
rect 30288 24896 30340 24948
rect 30564 24896 30616 24948
rect 34796 24939 34848 24948
rect 7748 24871 7800 24880
rect 7748 24837 7757 24871
rect 7757 24837 7791 24871
rect 7791 24837 7800 24871
rect 7748 24828 7800 24837
rect 8484 24828 8536 24880
rect 9680 24828 9732 24880
rect 10140 24828 10192 24880
rect 14740 24828 14792 24880
rect 19064 24871 19116 24880
rect 9956 24760 10008 24812
rect 11336 24760 11388 24812
rect 9588 24692 9640 24744
rect 12164 24735 12216 24744
rect 12164 24701 12173 24735
rect 12173 24701 12207 24735
rect 12207 24701 12216 24735
rect 12164 24692 12216 24701
rect 15292 24760 15344 24812
rect 19064 24837 19073 24871
rect 19073 24837 19107 24871
rect 19107 24837 19116 24871
rect 19064 24828 19116 24837
rect 20996 24871 21048 24880
rect 20996 24837 21005 24871
rect 21005 24837 21039 24871
rect 21039 24837 21048 24871
rect 20996 24828 21048 24837
rect 22284 24871 22336 24880
rect 22284 24837 22293 24871
rect 22293 24837 22327 24871
rect 22327 24837 22336 24871
rect 22284 24828 22336 24837
rect 25872 24828 25924 24880
rect 29092 24871 29144 24880
rect 29092 24837 29101 24871
rect 29101 24837 29135 24871
rect 29135 24837 29144 24871
rect 29092 24828 29144 24837
rect 12992 24735 13044 24744
rect 12992 24701 13001 24735
rect 13001 24701 13035 24735
rect 13035 24701 13044 24735
rect 12992 24692 13044 24701
rect 13176 24735 13228 24744
rect 13176 24701 13185 24735
rect 13185 24701 13219 24735
rect 13219 24701 13228 24735
rect 13176 24692 13228 24701
rect 15200 24692 15252 24744
rect 16764 24692 16816 24744
rect 9864 24624 9916 24676
rect 10876 24624 10928 24676
rect 10968 24624 11020 24676
rect 14464 24624 14516 24676
rect 9128 24556 9180 24608
rect 9220 24599 9272 24608
rect 9220 24565 9229 24599
rect 9229 24565 9263 24599
rect 9263 24565 9272 24599
rect 9220 24556 9272 24565
rect 10784 24556 10836 24608
rect 13544 24556 13596 24608
rect 17132 24556 17184 24608
rect 17868 24760 17920 24812
rect 19800 24760 19852 24812
rect 20352 24760 20404 24812
rect 23664 24760 23716 24812
rect 25780 24760 25832 24812
rect 27068 24760 27120 24812
rect 27436 24760 27488 24812
rect 27896 24803 27948 24812
rect 27896 24769 27905 24803
rect 27905 24769 27939 24803
rect 27939 24769 27948 24803
rect 27896 24760 27948 24769
rect 30748 24828 30800 24880
rect 31484 24828 31536 24880
rect 34796 24905 34805 24939
rect 34805 24905 34839 24939
rect 34839 24905 34848 24939
rect 34796 24896 34848 24905
rect 29736 24803 29788 24812
rect 29736 24769 29745 24803
rect 29745 24769 29779 24803
rect 29779 24769 29788 24803
rect 29736 24760 29788 24769
rect 30012 24760 30064 24812
rect 31208 24760 31260 24812
rect 18052 24692 18104 24744
rect 18236 24692 18288 24744
rect 18972 24692 19024 24744
rect 20812 24692 20864 24744
rect 21824 24692 21876 24744
rect 17960 24624 18012 24676
rect 18328 24556 18380 24608
rect 19984 24599 20036 24608
rect 19984 24565 19993 24599
rect 19993 24565 20027 24599
rect 20027 24565 20036 24599
rect 19984 24556 20036 24565
rect 22744 24556 22796 24608
rect 29460 24692 29512 24744
rect 29920 24692 29972 24744
rect 30656 24692 30708 24744
rect 32496 24760 32548 24812
rect 32220 24692 32272 24744
rect 33232 24760 33284 24812
rect 36360 24803 36412 24812
rect 33508 24692 33560 24744
rect 34704 24735 34756 24744
rect 27160 24556 27212 24608
rect 30472 24624 30524 24676
rect 31392 24624 31444 24676
rect 34704 24701 34713 24735
rect 34713 24701 34747 24735
rect 34747 24701 34756 24735
rect 34704 24692 34756 24701
rect 29000 24556 29052 24608
rect 29828 24556 29880 24608
rect 30012 24556 30064 24608
rect 30380 24556 30432 24608
rect 33784 24556 33836 24608
rect 33968 24599 34020 24608
rect 33968 24565 33977 24599
rect 33977 24565 34011 24599
rect 34011 24565 34020 24599
rect 33968 24556 34020 24565
rect 34612 24624 34664 24676
rect 36360 24769 36369 24803
rect 36369 24769 36403 24803
rect 36403 24769 36412 24803
rect 36360 24760 36412 24769
rect 36452 24803 36504 24812
rect 36452 24769 36461 24803
rect 36461 24769 36495 24803
rect 36495 24769 36504 24803
rect 36452 24760 36504 24769
rect 35348 24556 35400 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 7932 24352 7984 24404
rect 15660 24395 15712 24404
rect 15660 24361 15669 24395
rect 15669 24361 15703 24395
rect 15703 24361 15712 24395
rect 15660 24352 15712 24361
rect 16948 24352 17000 24404
rect 20352 24395 20404 24404
rect 8116 24284 8168 24336
rect 8208 24216 8260 24268
rect 11336 24284 11388 24336
rect 9128 24216 9180 24268
rect 9772 24216 9824 24268
rect 11152 24216 11204 24268
rect 11704 24216 11756 24268
rect 12348 24216 12400 24268
rect 17132 24259 17184 24268
rect 17132 24225 17141 24259
rect 17141 24225 17175 24259
rect 17175 24225 17184 24259
rect 17132 24216 17184 24225
rect 20352 24361 20361 24395
rect 20361 24361 20395 24395
rect 20395 24361 20404 24395
rect 20352 24352 20404 24361
rect 23664 24395 23716 24404
rect 23664 24361 23673 24395
rect 23673 24361 23707 24395
rect 23707 24361 23716 24395
rect 23664 24352 23716 24361
rect 27068 24395 27120 24404
rect 27068 24361 27077 24395
rect 27077 24361 27111 24395
rect 27111 24361 27120 24395
rect 27068 24352 27120 24361
rect 17868 24284 17920 24336
rect 30472 24352 30524 24404
rect 2228 24148 2280 24200
rect 9864 24148 9916 24200
rect 11336 24191 11388 24200
rect 11336 24157 11345 24191
rect 11345 24157 11379 24191
rect 11379 24157 11388 24191
rect 11336 24148 11388 24157
rect 13544 24191 13596 24200
rect 13544 24157 13553 24191
rect 13553 24157 13587 24191
rect 13587 24157 13596 24191
rect 13544 24148 13596 24157
rect 14464 24191 14516 24200
rect 14464 24157 14473 24191
rect 14473 24157 14507 24191
rect 14507 24157 14516 24191
rect 14464 24148 14516 24157
rect 18328 24191 18380 24200
rect 9220 24080 9272 24132
rect 11980 24123 12032 24132
rect 11980 24089 11989 24123
rect 11989 24089 12023 24123
rect 12023 24089 12032 24123
rect 11980 24080 12032 24089
rect 18328 24157 18337 24191
rect 18337 24157 18371 24191
rect 18371 24157 18380 24191
rect 18328 24148 18380 24157
rect 19616 24216 19668 24268
rect 19800 24216 19852 24268
rect 18604 24148 18656 24200
rect 20720 24148 20772 24200
rect 21180 24148 21232 24200
rect 1584 24055 1636 24064
rect 1584 24021 1593 24055
rect 1593 24021 1627 24055
rect 1627 24021 1636 24055
rect 1584 24012 1636 24021
rect 7288 24055 7340 24064
rect 7288 24021 7297 24055
rect 7297 24021 7331 24055
rect 7331 24021 7340 24055
rect 7288 24012 7340 24021
rect 11888 24012 11940 24064
rect 13268 24012 13320 24064
rect 14372 24055 14424 24064
rect 14372 24021 14381 24055
rect 14381 24021 14415 24055
rect 14415 24021 14424 24055
rect 14372 24012 14424 24021
rect 15476 24012 15528 24064
rect 16672 24080 16724 24132
rect 20904 24080 20956 24132
rect 25596 24216 25648 24268
rect 25872 24216 25924 24268
rect 26240 24216 26292 24268
rect 23112 24191 23164 24200
rect 23112 24157 23121 24191
rect 23121 24157 23155 24191
rect 23155 24157 23164 24191
rect 23112 24148 23164 24157
rect 24492 24148 24544 24200
rect 25504 24191 25556 24200
rect 25504 24157 25513 24191
rect 25513 24157 25547 24191
rect 25547 24157 25556 24191
rect 25504 24148 25556 24157
rect 28356 24148 28408 24200
rect 33508 24284 33560 24336
rect 30472 24216 30524 24268
rect 31944 24216 31996 24268
rect 32036 24216 32088 24268
rect 32312 24259 32364 24268
rect 32312 24225 32321 24259
rect 32321 24225 32355 24259
rect 32355 24225 32364 24259
rect 32312 24216 32364 24225
rect 32496 24216 32548 24268
rect 34704 24284 34756 24336
rect 34152 24259 34204 24268
rect 34152 24225 34161 24259
rect 34161 24225 34195 24259
rect 34195 24225 34204 24259
rect 34152 24216 34204 24225
rect 34612 24216 34664 24268
rect 32220 24148 32272 24200
rect 33140 24148 33192 24200
rect 36912 24191 36964 24200
rect 36912 24157 36921 24191
rect 36921 24157 36955 24191
rect 36955 24157 36964 24191
rect 36912 24148 36964 24157
rect 36820 24080 36872 24132
rect 17776 24012 17828 24064
rect 19892 24012 19944 24064
rect 21088 24012 21140 24064
rect 22560 24012 22612 24064
rect 24400 24012 24452 24064
rect 26148 24012 26200 24064
rect 33600 24012 33652 24064
rect 34428 24012 34480 24064
rect 34980 24012 35032 24064
rect 37096 24055 37148 24064
rect 37096 24021 37105 24055
rect 37105 24021 37139 24055
rect 37139 24021 37148 24055
rect 37096 24012 37148 24021
rect 4874 23910 4926 23962
rect 4938 23910 4990 23962
rect 5002 23910 5054 23962
rect 5066 23910 5118 23962
rect 5130 23910 5182 23962
rect 35594 23910 35646 23962
rect 35658 23910 35710 23962
rect 35722 23910 35774 23962
rect 35786 23910 35838 23962
rect 35850 23910 35902 23962
rect 9312 23808 9364 23860
rect 10784 23851 10836 23860
rect 10784 23817 10793 23851
rect 10793 23817 10827 23851
rect 10827 23817 10836 23851
rect 10784 23808 10836 23817
rect 12164 23851 12216 23860
rect 12164 23817 12173 23851
rect 12173 23817 12207 23851
rect 12207 23817 12216 23851
rect 12164 23808 12216 23817
rect 14740 23851 14792 23860
rect 7288 23740 7340 23792
rect 10232 23740 10284 23792
rect 14740 23817 14749 23851
rect 14749 23817 14783 23851
rect 14783 23817 14792 23851
rect 14740 23808 14792 23817
rect 16580 23808 16632 23860
rect 16672 23808 16724 23860
rect 13268 23783 13320 23792
rect 13268 23749 13277 23783
rect 13277 23749 13311 23783
rect 13311 23749 13320 23783
rect 13268 23740 13320 23749
rect 6920 23604 6972 23656
rect 7288 23647 7340 23656
rect 7288 23613 7297 23647
rect 7297 23613 7331 23647
rect 7331 23613 7340 23647
rect 7288 23604 7340 23613
rect 8760 23647 8812 23656
rect 8760 23613 8769 23647
rect 8769 23613 8803 23647
rect 8803 23613 8812 23647
rect 8760 23604 8812 23613
rect 9680 23647 9732 23656
rect 9680 23613 9689 23647
rect 9689 23613 9723 23647
rect 9723 23613 9732 23647
rect 9680 23604 9732 23613
rect 9772 23647 9824 23656
rect 9772 23613 9781 23647
rect 9781 23613 9815 23647
rect 9815 23613 9824 23647
rect 9772 23604 9824 23613
rect 11796 23604 11848 23656
rect 12348 23672 12400 23724
rect 14372 23672 14424 23724
rect 15200 23672 15252 23724
rect 16764 23672 16816 23724
rect 17868 23808 17920 23860
rect 19800 23808 19852 23860
rect 20812 23808 20864 23860
rect 17776 23783 17828 23792
rect 17776 23749 17785 23783
rect 17785 23749 17819 23783
rect 17819 23749 17828 23783
rect 17776 23740 17828 23749
rect 18512 23740 18564 23792
rect 19984 23783 20036 23792
rect 19984 23749 19993 23783
rect 19993 23749 20027 23783
rect 20027 23749 20036 23783
rect 19984 23740 20036 23749
rect 21088 23672 21140 23724
rect 23112 23808 23164 23860
rect 24400 23851 24452 23860
rect 24400 23817 24409 23851
rect 24409 23817 24443 23851
rect 24443 23817 24452 23851
rect 24400 23808 24452 23817
rect 26148 23851 26200 23860
rect 26148 23817 26157 23851
rect 26157 23817 26191 23851
rect 26191 23817 26200 23851
rect 26148 23808 26200 23817
rect 28080 23808 28132 23860
rect 33232 23808 33284 23860
rect 36820 23851 36872 23860
rect 36820 23817 36829 23851
rect 36829 23817 36863 23851
rect 36863 23817 36872 23851
rect 36820 23808 36872 23817
rect 27896 23740 27948 23792
rect 30472 23740 30524 23792
rect 22836 23715 22888 23724
rect 22836 23681 22845 23715
rect 22845 23681 22879 23715
rect 22879 23681 22888 23715
rect 22836 23672 22888 23681
rect 32496 23715 32548 23724
rect 9588 23536 9640 23588
rect 14004 23604 14056 23656
rect 19708 23647 19760 23656
rect 12348 23536 12400 23588
rect 9312 23468 9364 23520
rect 10600 23468 10652 23520
rect 12532 23511 12584 23520
rect 12532 23477 12541 23511
rect 12541 23477 12575 23511
rect 12575 23477 12584 23511
rect 12532 23468 12584 23477
rect 19708 23613 19717 23647
rect 19717 23613 19751 23647
rect 19751 23613 19760 23647
rect 19708 23604 19760 23613
rect 23848 23604 23900 23656
rect 24676 23647 24728 23656
rect 24676 23613 24685 23647
rect 24685 23613 24719 23647
rect 24719 23613 24728 23647
rect 24676 23604 24728 23613
rect 25688 23604 25740 23656
rect 25872 23647 25924 23656
rect 25872 23613 25881 23647
rect 25881 23613 25915 23647
rect 25915 23613 25924 23647
rect 25872 23604 25924 23613
rect 26056 23647 26108 23656
rect 26056 23613 26065 23647
rect 26065 23613 26099 23647
rect 26099 23613 26108 23647
rect 26056 23604 26108 23613
rect 27160 23647 27212 23656
rect 27160 23613 27169 23647
rect 27169 23613 27203 23647
rect 27203 23613 27212 23647
rect 27160 23604 27212 23613
rect 27436 23647 27488 23656
rect 27436 23613 27445 23647
rect 27445 23613 27479 23647
rect 27479 23613 27488 23647
rect 27436 23604 27488 23613
rect 30104 23647 30156 23656
rect 30104 23613 30113 23647
rect 30113 23613 30147 23647
rect 30147 23613 30156 23647
rect 30104 23604 30156 23613
rect 32496 23681 32505 23715
rect 32505 23681 32539 23715
rect 32539 23681 32548 23715
rect 32496 23672 32548 23681
rect 33508 23715 33560 23724
rect 33508 23681 33517 23715
rect 33517 23681 33551 23715
rect 33551 23681 33560 23715
rect 33508 23672 33560 23681
rect 34428 23715 34480 23724
rect 34428 23681 34437 23715
rect 34437 23681 34471 23715
rect 34471 23681 34480 23715
rect 34428 23672 34480 23681
rect 31944 23604 31996 23656
rect 32404 23647 32456 23656
rect 32404 23613 32413 23647
rect 32413 23613 32447 23647
rect 32447 23613 32456 23647
rect 32404 23604 32456 23613
rect 33600 23647 33652 23656
rect 33600 23613 33609 23647
rect 33609 23613 33643 23647
rect 33643 23613 33652 23647
rect 33600 23604 33652 23613
rect 34980 23672 35032 23724
rect 35440 23740 35492 23792
rect 36452 23672 36504 23724
rect 16212 23468 16264 23520
rect 20168 23468 20220 23520
rect 21456 23511 21508 23520
rect 21456 23477 21465 23511
rect 21465 23477 21499 23511
rect 21499 23477 21508 23511
rect 21456 23468 21508 23477
rect 26332 23468 26384 23520
rect 32128 23468 32180 23520
rect 32312 23468 32364 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 7288 23264 7340 23316
rect 7564 23264 7616 23316
rect 11336 23264 11388 23316
rect 13912 23264 13964 23316
rect 18512 23264 18564 23316
rect 19064 23264 19116 23316
rect 19616 23264 19668 23316
rect 20260 23264 20312 23316
rect 20996 23264 21048 23316
rect 9772 23196 9824 23248
rect 12164 23196 12216 23248
rect 12440 23196 12492 23248
rect 13084 23196 13136 23248
rect 27436 23264 27488 23316
rect 27896 23264 27948 23316
rect 29092 23264 29144 23316
rect 30472 23307 30524 23316
rect 30472 23273 30481 23307
rect 30481 23273 30515 23307
rect 30515 23273 30524 23307
rect 30472 23264 30524 23273
rect 31944 23264 31996 23316
rect 32772 23264 32824 23316
rect 33508 23264 33560 23316
rect 34704 23264 34756 23316
rect 8116 23128 8168 23180
rect 9588 23128 9640 23180
rect 11520 23128 11572 23180
rect 11796 23128 11848 23180
rect 13176 23171 13228 23180
rect 7564 22992 7616 23044
rect 6920 22967 6972 22976
rect 6920 22933 6929 22967
rect 6929 22933 6963 22967
rect 6963 22933 6972 22967
rect 6920 22924 6972 22933
rect 7472 22924 7524 22976
rect 8576 23060 8628 23112
rect 10784 23035 10836 23044
rect 10784 23001 10793 23035
rect 10793 23001 10827 23035
rect 10827 23001 10836 23035
rect 10784 22992 10836 23001
rect 12072 22992 12124 23044
rect 13176 23137 13185 23171
rect 13185 23137 13219 23171
rect 13219 23137 13228 23171
rect 13176 23128 13228 23137
rect 12532 23060 12584 23112
rect 12624 22992 12676 23044
rect 15476 23128 15528 23180
rect 17592 23128 17644 23180
rect 19892 23128 19944 23180
rect 16764 23103 16816 23112
rect 16764 23069 16773 23103
rect 16773 23069 16807 23103
rect 16807 23069 16816 23103
rect 16764 23060 16816 23069
rect 17500 23060 17552 23112
rect 17960 23060 18012 23112
rect 19248 23060 19300 23112
rect 20168 23171 20220 23180
rect 20168 23137 20177 23171
rect 20177 23137 20211 23171
rect 20211 23137 20220 23171
rect 20168 23128 20220 23137
rect 20996 23128 21048 23180
rect 21824 23128 21876 23180
rect 22652 23128 22704 23180
rect 25596 23171 25648 23180
rect 21456 23103 21508 23112
rect 21456 23069 21465 23103
rect 21465 23069 21499 23103
rect 21499 23069 21508 23103
rect 21456 23060 21508 23069
rect 25596 23137 25605 23171
rect 25605 23137 25639 23171
rect 25639 23137 25648 23171
rect 25596 23128 25648 23137
rect 26056 23060 26108 23112
rect 26332 23103 26384 23112
rect 26332 23069 26341 23103
rect 26341 23069 26375 23103
rect 26375 23069 26384 23103
rect 26332 23060 26384 23069
rect 27712 23103 27764 23112
rect 27712 23069 27721 23103
rect 27721 23069 27755 23103
rect 27755 23069 27764 23103
rect 27712 23060 27764 23069
rect 8760 22924 8812 22976
rect 9220 22924 9272 22976
rect 13912 22924 13964 22976
rect 22560 23035 22612 23044
rect 17316 22967 17368 22976
rect 17316 22933 17325 22967
rect 17325 22933 17359 22967
rect 17359 22933 17368 22967
rect 17316 22924 17368 22933
rect 19892 22967 19944 22976
rect 19892 22933 19901 22967
rect 19901 22933 19935 22967
rect 19935 22933 19944 22967
rect 19892 22924 19944 22933
rect 20904 22924 20956 22976
rect 22560 23001 22569 23035
rect 22569 23001 22603 23035
rect 22603 23001 22612 23035
rect 22560 22992 22612 23001
rect 23572 22992 23624 23044
rect 29736 23103 29788 23112
rect 28448 23035 28500 23044
rect 28448 23001 28457 23035
rect 28457 23001 28491 23035
rect 28491 23001 28500 23035
rect 28448 22992 28500 23001
rect 29736 23069 29745 23103
rect 29745 23069 29779 23103
rect 29779 23069 29788 23103
rect 29736 23060 29788 23069
rect 30564 23060 30616 23112
rect 30656 22992 30708 23044
rect 32496 23128 32548 23180
rect 35440 23128 35492 23180
rect 33600 23103 33652 23112
rect 33600 23069 33609 23103
rect 33609 23069 33643 23103
rect 33643 23069 33652 23103
rect 33600 23060 33652 23069
rect 33784 23103 33836 23112
rect 33784 23069 33793 23103
rect 33793 23069 33827 23103
rect 33827 23069 33836 23103
rect 33784 23060 33836 23069
rect 32220 22992 32272 23044
rect 32956 23035 33008 23044
rect 32956 23001 32965 23035
rect 32965 23001 32999 23035
rect 32999 23001 33008 23035
rect 32956 22992 33008 23001
rect 35348 22992 35400 23044
rect 25320 22924 25372 22976
rect 25964 22924 26016 22976
rect 27988 22924 28040 22976
rect 28632 22967 28684 22976
rect 28632 22933 28641 22967
rect 28641 22933 28675 22967
rect 28675 22933 28684 22967
rect 28632 22924 28684 22933
rect 29828 22967 29880 22976
rect 29828 22933 29837 22967
rect 29837 22933 29871 22967
rect 29871 22933 29880 22967
rect 29828 22924 29880 22933
rect 30564 22924 30616 22976
rect 31116 22924 31168 22976
rect 35992 22924 36044 22976
rect 4874 22822 4926 22874
rect 4938 22822 4990 22874
rect 5002 22822 5054 22874
rect 5066 22822 5118 22874
rect 5130 22822 5182 22874
rect 35594 22822 35646 22874
rect 35658 22822 35710 22874
rect 35722 22822 35774 22874
rect 35786 22822 35838 22874
rect 35850 22822 35902 22874
rect 6920 22720 6972 22772
rect 8208 22720 8260 22772
rect 9680 22720 9732 22772
rect 13268 22720 13320 22772
rect 6828 22652 6880 22704
rect 10048 22652 10100 22704
rect 11888 22652 11940 22704
rect 12440 22652 12492 22704
rect 14648 22652 14700 22704
rect 14924 22695 14976 22704
rect 14924 22661 14933 22695
rect 14933 22661 14967 22695
rect 14967 22661 14976 22695
rect 14924 22652 14976 22661
rect 8024 22584 8076 22636
rect 9128 22627 9180 22636
rect 9128 22593 9137 22627
rect 9137 22593 9171 22627
rect 9171 22593 9180 22627
rect 9128 22584 9180 22593
rect 11704 22627 11756 22636
rect 11704 22593 11713 22627
rect 11713 22593 11747 22627
rect 11747 22593 11756 22627
rect 11704 22584 11756 22593
rect 13912 22627 13964 22636
rect 13912 22593 13921 22627
rect 13921 22593 13955 22627
rect 13955 22593 13964 22627
rect 13912 22584 13964 22593
rect 21916 22720 21968 22772
rect 25320 22763 25372 22772
rect 25320 22729 25329 22763
rect 25329 22729 25363 22763
rect 25363 22729 25372 22763
rect 25320 22720 25372 22729
rect 17316 22652 17368 22704
rect 23664 22652 23716 22704
rect 28080 22720 28132 22772
rect 27896 22652 27948 22704
rect 18604 22627 18656 22636
rect 18604 22593 18613 22627
rect 18613 22593 18647 22627
rect 18647 22593 18656 22627
rect 18604 22584 18656 22593
rect 19248 22584 19300 22636
rect 20536 22627 20588 22636
rect 20536 22593 20545 22627
rect 20545 22593 20579 22627
rect 20579 22593 20588 22627
rect 20536 22584 20588 22593
rect 21180 22584 21232 22636
rect 22744 22627 22796 22636
rect 22744 22593 22753 22627
rect 22753 22593 22787 22627
rect 22787 22593 22796 22627
rect 22744 22584 22796 22593
rect 24676 22584 24728 22636
rect 26148 22627 26200 22636
rect 6920 22559 6972 22568
rect 6920 22525 6929 22559
rect 6929 22525 6963 22559
rect 6963 22525 6972 22559
rect 9404 22559 9456 22568
rect 6920 22516 6972 22525
rect 9404 22525 9413 22559
rect 9413 22525 9447 22559
rect 9447 22525 9456 22559
rect 9404 22516 9456 22525
rect 14004 22448 14056 22500
rect 14096 22423 14148 22432
rect 14096 22389 14105 22423
rect 14105 22389 14139 22423
rect 14139 22389 14148 22423
rect 14096 22380 14148 22389
rect 15568 22448 15620 22500
rect 19892 22516 19944 22568
rect 23020 22559 23072 22568
rect 20260 22448 20312 22500
rect 23020 22525 23029 22559
rect 23029 22525 23063 22559
rect 23063 22525 23072 22559
rect 23020 22516 23072 22525
rect 25412 22559 25464 22568
rect 25412 22525 25421 22559
rect 25421 22525 25455 22559
rect 25455 22525 25464 22559
rect 25412 22516 25464 22525
rect 26148 22593 26157 22627
rect 26157 22593 26191 22627
rect 26191 22593 26200 22627
rect 26148 22584 26200 22593
rect 33140 22720 33192 22772
rect 35992 22720 36044 22772
rect 36452 22763 36504 22772
rect 36452 22729 36461 22763
rect 36461 22729 36495 22763
rect 36495 22729 36504 22763
rect 36452 22720 36504 22729
rect 30656 22695 30708 22704
rect 30656 22661 30665 22695
rect 30665 22661 30699 22695
rect 30699 22661 30708 22695
rect 30656 22652 30708 22661
rect 31760 22652 31812 22704
rect 32772 22695 32824 22704
rect 32772 22661 32807 22695
rect 32807 22661 32824 22695
rect 32772 22652 32824 22661
rect 32956 22652 33008 22704
rect 36084 22652 36136 22704
rect 30748 22627 30800 22636
rect 30748 22593 30757 22627
rect 30757 22593 30791 22627
rect 30791 22593 30800 22627
rect 30748 22584 30800 22593
rect 27160 22559 27212 22568
rect 27160 22525 27169 22559
rect 27169 22525 27203 22559
rect 27203 22525 27212 22559
rect 27160 22516 27212 22525
rect 30380 22448 30432 22500
rect 33692 22584 33744 22636
rect 36544 22627 36596 22636
rect 36544 22593 36553 22627
rect 36553 22593 36587 22627
rect 36587 22593 36596 22627
rect 36544 22584 36596 22593
rect 33140 22516 33192 22568
rect 35256 22516 35308 22568
rect 17592 22380 17644 22432
rect 18604 22380 18656 22432
rect 19248 22423 19300 22432
rect 19248 22389 19257 22423
rect 19257 22389 19291 22423
rect 19291 22389 19300 22423
rect 19248 22380 19300 22389
rect 20168 22423 20220 22432
rect 20168 22389 20177 22423
rect 20177 22389 20211 22423
rect 20211 22389 20220 22423
rect 20168 22380 20220 22389
rect 22100 22423 22152 22432
rect 22100 22389 22109 22423
rect 22109 22389 22143 22423
rect 22143 22389 22152 22423
rect 24952 22423 25004 22432
rect 22100 22380 22152 22389
rect 24952 22389 24961 22423
rect 24961 22389 24995 22423
rect 24995 22389 25004 22423
rect 24952 22380 25004 22389
rect 29736 22423 29788 22432
rect 29736 22389 29745 22423
rect 29745 22389 29779 22423
rect 29779 22389 29788 22423
rect 29736 22380 29788 22389
rect 33968 22448 34020 22500
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 6920 22176 6972 22228
rect 9404 22176 9456 22228
rect 10784 22219 10836 22228
rect 10784 22185 10793 22219
rect 10793 22185 10827 22219
rect 10827 22185 10836 22219
rect 10784 22176 10836 22185
rect 14096 22176 14148 22228
rect 17684 22176 17736 22228
rect 20260 22176 20312 22228
rect 31944 22219 31996 22228
rect 31944 22185 31953 22219
rect 31953 22185 31987 22219
rect 31987 22185 31996 22219
rect 31944 22176 31996 22185
rect 32588 22176 32640 22228
rect 33508 22176 33560 22228
rect 34428 22176 34480 22228
rect 11704 22108 11756 22160
rect 8024 22083 8076 22092
rect 8024 22049 8033 22083
rect 8033 22049 8067 22083
rect 8067 22049 8076 22083
rect 8024 22040 8076 22049
rect 7472 22015 7524 22024
rect 7472 21981 7481 22015
rect 7481 21981 7515 22015
rect 7515 21981 7524 22015
rect 7472 21972 7524 21981
rect 8300 22040 8352 22092
rect 10048 22083 10100 22092
rect 10048 22049 10057 22083
rect 10057 22049 10091 22083
rect 10091 22049 10100 22083
rect 10048 22040 10100 22049
rect 12440 22040 12492 22092
rect 13084 22083 13136 22092
rect 13084 22049 13093 22083
rect 13093 22049 13127 22083
rect 13127 22049 13136 22083
rect 13084 22040 13136 22049
rect 15568 22108 15620 22160
rect 9312 22015 9364 22024
rect 9312 21981 9321 22015
rect 9321 21981 9355 22015
rect 9355 21981 9364 22015
rect 9312 21972 9364 21981
rect 9496 21972 9548 22024
rect 10600 22015 10652 22024
rect 10600 21981 10609 22015
rect 10609 21981 10643 22015
rect 10643 21981 10652 22015
rect 10600 21972 10652 21981
rect 12164 21972 12216 22024
rect 13176 21972 13228 22024
rect 14924 22040 14976 22092
rect 14096 21972 14148 22024
rect 15016 21904 15068 21956
rect 17684 22040 17736 22092
rect 18972 22108 19024 22160
rect 17500 21972 17552 22024
rect 18236 21972 18288 22024
rect 19892 22108 19944 22160
rect 28448 22108 28500 22160
rect 19800 22040 19852 22092
rect 23572 22040 23624 22092
rect 20168 21972 20220 22024
rect 22100 21972 22152 22024
rect 24952 22040 25004 22092
rect 25688 22083 25740 22092
rect 25688 22049 25697 22083
rect 25697 22049 25731 22083
rect 25731 22049 25740 22083
rect 25688 22040 25740 22049
rect 27896 22040 27948 22092
rect 28724 22083 28776 22092
rect 28724 22049 28733 22083
rect 28733 22049 28767 22083
rect 28767 22049 28776 22083
rect 28724 22040 28776 22049
rect 30288 22083 30340 22092
rect 17132 21904 17184 21956
rect 12440 21836 12492 21888
rect 12808 21836 12860 21888
rect 12992 21879 13044 21888
rect 12992 21845 13001 21879
rect 13001 21845 13035 21879
rect 13035 21845 13044 21879
rect 12992 21836 13044 21845
rect 16028 21879 16080 21888
rect 16028 21845 16037 21879
rect 16037 21845 16071 21879
rect 16071 21845 16080 21879
rect 16028 21836 16080 21845
rect 16672 21879 16724 21888
rect 16672 21845 16681 21879
rect 16681 21845 16715 21879
rect 16715 21845 16724 21879
rect 16672 21836 16724 21845
rect 18696 21836 18748 21888
rect 18880 21879 18932 21888
rect 18880 21845 18889 21879
rect 18889 21845 18923 21879
rect 18923 21845 18932 21879
rect 18880 21836 18932 21845
rect 24492 21972 24544 22024
rect 25964 22015 26016 22024
rect 25964 21981 25973 22015
rect 25973 21981 26007 22015
rect 26007 21981 26016 22015
rect 25964 21972 26016 21981
rect 27712 21972 27764 22024
rect 29368 21972 29420 22024
rect 29552 21972 29604 22024
rect 29828 21972 29880 22024
rect 30288 22049 30297 22083
rect 30297 22049 30331 22083
rect 30331 22049 30340 22083
rect 30288 22040 30340 22049
rect 31760 22040 31812 22092
rect 30380 21972 30432 22024
rect 23572 21904 23624 21956
rect 25412 21904 25464 21956
rect 31944 21972 31996 22024
rect 33600 22108 33652 22160
rect 34796 22108 34848 22160
rect 32404 22040 32456 22092
rect 33692 22040 33744 22092
rect 33600 22015 33652 22024
rect 33600 21981 33609 22015
rect 33609 21981 33643 22015
rect 33643 21981 33652 22015
rect 33600 21972 33652 21981
rect 34428 22040 34480 22092
rect 35348 22040 35400 22092
rect 33968 22015 34020 22024
rect 33968 21981 33977 22015
rect 33977 21981 34011 22015
rect 34011 21981 34020 22015
rect 33968 21972 34020 21981
rect 32864 21904 32916 21956
rect 33140 21904 33192 21956
rect 36084 21972 36136 22024
rect 36544 21972 36596 22024
rect 22008 21836 22060 21888
rect 23020 21836 23072 21888
rect 24676 21879 24728 21888
rect 24676 21845 24685 21879
rect 24685 21845 24719 21879
rect 24719 21845 24728 21879
rect 24676 21836 24728 21845
rect 26148 21836 26200 21888
rect 26976 21879 27028 21888
rect 26976 21845 26985 21879
rect 26985 21845 27019 21879
rect 27019 21845 27028 21879
rect 26976 21836 27028 21845
rect 29184 21879 29236 21888
rect 29184 21845 29193 21879
rect 29193 21845 29227 21879
rect 29227 21845 29236 21879
rect 29184 21836 29236 21845
rect 33416 21879 33468 21888
rect 33416 21845 33425 21879
rect 33425 21845 33459 21879
rect 33459 21845 33468 21879
rect 33416 21836 33468 21845
rect 33600 21836 33652 21888
rect 35992 21836 36044 21888
rect 4874 21734 4926 21786
rect 4938 21734 4990 21786
rect 5002 21734 5054 21786
rect 5066 21734 5118 21786
rect 5130 21734 5182 21786
rect 35594 21734 35646 21786
rect 35658 21734 35710 21786
rect 35722 21734 35774 21786
rect 35786 21734 35838 21786
rect 35850 21734 35902 21786
rect 12072 21675 12124 21684
rect 12072 21641 12081 21675
rect 12081 21641 12115 21675
rect 12115 21641 12124 21675
rect 12072 21632 12124 21641
rect 13912 21675 13964 21684
rect 13912 21641 13921 21675
rect 13921 21641 13955 21675
rect 13955 21641 13964 21675
rect 13912 21632 13964 21641
rect 15016 21632 15068 21684
rect 18236 21675 18288 21684
rect 18236 21641 18245 21675
rect 18245 21641 18279 21675
rect 18279 21641 18288 21675
rect 18236 21632 18288 21641
rect 18696 21632 18748 21684
rect 20536 21632 20588 21684
rect 22008 21632 22060 21684
rect 23664 21675 23716 21684
rect 23664 21641 23673 21675
rect 23673 21641 23707 21675
rect 23707 21641 23716 21675
rect 23664 21632 23716 21641
rect 25412 21632 25464 21684
rect 27252 21632 27304 21684
rect 29552 21675 29604 21684
rect 29552 21641 29561 21675
rect 29561 21641 29595 21675
rect 29595 21641 29604 21675
rect 29552 21632 29604 21641
rect 30288 21632 30340 21684
rect 32864 21675 32916 21684
rect 32864 21641 32873 21675
rect 32873 21641 32907 21675
rect 32907 21641 32916 21675
rect 32864 21632 32916 21641
rect 12992 21564 13044 21616
rect 16028 21564 16080 21616
rect 17500 21564 17552 21616
rect 19248 21564 19300 21616
rect 19800 21564 19852 21616
rect 8300 21496 8352 21548
rect 10140 21539 10192 21548
rect 10140 21505 10149 21539
rect 10149 21505 10183 21539
rect 10183 21505 10192 21539
rect 10140 21496 10192 21505
rect 12164 21539 12216 21548
rect 12164 21505 12173 21539
rect 12173 21505 12207 21539
rect 12207 21505 12216 21539
rect 12164 21496 12216 21505
rect 14372 21496 14424 21548
rect 15844 21539 15896 21548
rect 15844 21505 15853 21539
rect 15853 21505 15887 21539
rect 15887 21505 15896 21539
rect 15844 21496 15896 21505
rect 17776 21496 17828 21548
rect 26976 21564 27028 21616
rect 29736 21564 29788 21616
rect 21088 21496 21140 21548
rect 23572 21539 23624 21548
rect 13268 21471 13320 21480
rect 13268 21437 13277 21471
rect 13277 21437 13311 21471
rect 13311 21437 13320 21471
rect 13268 21428 13320 21437
rect 13452 21471 13504 21480
rect 13452 21437 13461 21471
rect 13461 21437 13495 21471
rect 13495 21437 13504 21471
rect 13452 21428 13504 21437
rect 16488 21428 16540 21480
rect 17960 21428 18012 21480
rect 18236 21428 18288 21480
rect 19708 21471 19760 21480
rect 19708 21437 19717 21471
rect 19717 21437 19751 21471
rect 19751 21437 19760 21471
rect 19708 21428 19760 21437
rect 20996 21471 21048 21480
rect 20996 21437 21005 21471
rect 21005 21437 21039 21471
rect 21039 21437 21048 21471
rect 20996 21428 21048 21437
rect 21824 21428 21876 21480
rect 14740 21360 14792 21412
rect 21916 21360 21968 21412
rect 23572 21505 23581 21539
rect 23581 21505 23615 21539
rect 23615 21505 23624 21539
rect 23572 21496 23624 21505
rect 24492 21496 24544 21548
rect 26516 21496 26568 21548
rect 27160 21539 27212 21548
rect 27160 21505 27169 21539
rect 27169 21505 27203 21539
rect 27203 21505 27212 21539
rect 27160 21496 27212 21505
rect 30380 21564 30432 21616
rect 33508 21564 33560 21616
rect 35992 21564 36044 21616
rect 25596 21428 25648 21480
rect 25780 21471 25832 21480
rect 25780 21437 25789 21471
rect 25789 21437 25823 21471
rect 25823 21437 25832 21471
rect 25780 21428 25832 21437
rect 30564 21496 30616 21548
rect 32496 21539 32548 21548
rect 7840 21292 7892 21344
rect 9956 21335 10008 21344
rect 9956 21301 9965 21335
rect 9965 21301 9999 21335
rect 9999 21301 10008 21335
rect 9956 21292 10008 21301
rect 16488 21292 16540 21344
rect 18696 21292 18748 21344
rect 24308 21335 24360 21344
rect 24308 21301 24317 21335
rect 24317 21301 24351 21335
rect 24351 21301 24360 21335
rect 24308 21292 24360 21301
rect 24952 21292 25004 21344
rect 29368 21403 29420 21412
rect 29368 21369 29377 21403
rect 29377 21369 29411 21403
rect 29411 21369 29420 21403
rect 29368 21360 29420 21369
rect 30472 21428 30524 21480
rect 32496 21505 32505 21539
rect 32505 21505 32539 21539
rect 32539 21505 32548 21539
rect 32496 21496 32548 21505
rect 32588 21496 32640 21548
rect 32404 21471 32456 21480
rect 32404 21437 32413 21471
rect 32413 21437 32447 21471
rect 32447 21437 32456 21471
rect 32404 21428 32456 21437
rect 33692 21471 33744 21480
rect 33692 21437 33701 21471
rect 33701 21437 33735 21471
rect 33735 21437 33744 21471
rect 33692 21428 33744 21437
rect 34336 21428 34388 21480
rect 35348 21428 35400 21480
rect 31484 21360 31536 21412
rect 28632 21292 28684 21344
rect 30288 21292 30340 21344
rect 30380 21292 30432 21344
rect 30840 21335 30892 21344
rect 30840 21301 30849 21335
rect 30849 21301 30883 21335
rect 30883 21301 30892 21335
rect 30840 21292 30892 21301
rect 34060 21335 34112 21344
rect 34060 21301 34069 21335
rect 34069 21301 34103 21335
rect 34103 21301 34112 21335
rect 34060 21292 34112 21301
rect 34796 21292 34848 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 8576 21131 8628 21140
rect 8576 21097 8585 21131
rect 8585 21097 8619 21131
rect 8619 21097 8628 21131
rect 8576 21088 8628 21097
rect 15844 21088 15896 21140
rect 26516 21131 26568 21140
rect 9588 21020 9640 21072
rect 11980 21020 12032 21072
rect 12532 21020 12584 21072
rect 26516 21097 26525 21131
rect 26525 21097 26559 21131
rect 26559 21097 26568 21131
rect 26516 21088 26568 21097
rect 28724 21131 28776 21140
rect 28724 21097 28733 21131
rect 28733 21097 28767 21131
rect 28767 21097 28776 21131
rect 28724 21088 28776 21097
rect 6828 20995 6880 21004
rect 6828 20961 6837 20995
rect 6837 20961 6871 20995
rect 6871 20961 6880 20995
rect 6828 20952 6880 20961
rect 10876 20952 10928 21004
rect 12624 20995 12676 21004
rect 9588 20884 9640 20936
rect 7104 20859 7156 20868
rect 7104 20825 7113 20859
rect 7113 20825 7147 20859
rect 7147 20825 7156 20859
rect 7104 20816 7156 20825
rect 7840 20816 7892 20868
rect 8760 20816 8812 20868
rect 8668 20748 8720 20800
rect 10784 20748 10836 20800
rect 11612 20791 11664 20800
rect 11612 20757 11621 20791
rect 11621 20757 11655 20791
rect 11655 20757 11664 20791
rect 11612 20748 11664 20757
rect 12624 20961 12633 20995
rect 12633 20961 12667 20995
rect 12667 20961 12676 20995
rect 12624 20952 12676 20961
rect 26792 21020 26844 21072
rect 20076 20952 20128 21004
rect 20720 20952 20772 21004
rect 21824 20952 21876 21004
rect 23572 20952 23624 21004
rect 25136 20995 25188 21004
rect 25136 20961 25145 20995
rect 25145 20961 25179 20995
rect 25179 20961 25188 20995
rect 25136 20952 25188 20961
rect 25320 20952 25372 21004
rect 25688 20952 25740 21004
rect 12440 20927 12492 20936
rect 12440 20893 12449 20927
rect 12449 20893 12483 20927
rect 12483 20893 12492 20927
rect 14280 20927 14332 20936
rect 12440 20884 12492 20893
rect 14280 20893 14289 20927
rect 14289 20893 14323 20927
rect 14323 20893 14332 20927
rect 14280 20884 14332 20893
rect 14372 20884 14424 20936
rect 17684 20927 17736 20936
rect 17684 20893 17693 20927
rect 17693 20893 17727 20927
rect 17727 20893 17736 20927
rect 17684 20884 17736 20893
rect 19892 20884 19944 20936
rect 24952 20927 25004 20936
rect 24952 20893 24961 20927
rect 24961 20893 24995 20927
rect 24995 20893 25004 20927
rect 24952 20884 25004 20893
rect 27528 20952 27580 21004
rect 32404 21088 32456 21140
rect 33692 21088 33744 21140
rect 31484 21020 31536 21072
rect 31208 20952 31260 21004
rect 34612 21020 34664 21072
rect 34796 20952 34848 21004
rect 16672 20816 16724 20868
rect 17408 20859 17460 20868
rect 17408 20825 17417 20859
rect 17417 20825 17451 20859
rect 17451 20825 17460 20859
rect 17408 20816 17460 20825
rect 18052 20816 18104 20868
rect 18512 20859 18564 20868
rect 18512 20825 18521 20859
rect 18521 20825 18555 20859
rect 18555 20825 18564 20859
rect 18512 20816 18564 20825
rect 21364 20859 21416 20868
rect 21364 20825 21373 20859
rect 21373 20825 21407 20859
rect 21407 20825 21416 20859
rect 21364 20816 21416 20825
rect 13452 20748 13504 20800
rect 14464 20791 14516 20800
rect 14464 20757 14473 20791
rect 14473 20757 14507 20791
rect 14507 20757 14516 20791
rect 14464 20748 14516 20757
rect 15384 20748 15436 20800
rect 15660 20748 15712 20800
rect 17776 20748 17828 20800
rect 22100 20816 22152 20868
rect 28448 20884 28500 20936
rect 29000 20927 29052 20936
rect 29000 20893 29009 20927
rect 29009 20893 29043 20927
rect 29043 20893 29052 20927
rect 29000 20884 29052 20893
rect 29736 20884 29788 20936
rect 31576 20884 31628 20936
rect 27712 20816 27764 20868
rect 28724 20816 28776 20868
rect 30472 20859 30524 20868
rect 30472 20825 30481 20859
rect 30481 20825 30515 20859
rect 30515 20825 30524 20859
rect 30472 20816 30524 20825
rect 32864 20884 32916 20936
rect 33600 20884 33652 20936
rect 34060 20884 34112 20936
rect 33416 20816 33468 20868
rect 33508 20816 33560 20868
rect 21824 20791 21876 20800
rect 21824 20757 21833 20791
rect 21833 20757 21867 20791
rect 21867 20757 21876 20791
rect 21824 20748 21876 20757
rect 22284 20791 22336 20800
rect 22284 20757 22293 20791
rect 22293 20757 22327 20791
rect 22327 20757 22336 20791
rect 22284 20748 22336 20757
rect 24768 20748 24820 20800
rect 25596 20748 25648 20800
rect 27252 20748 27304 20800
rect 30564 20748 30616 20800
rect 33784 20791 33836 20800
rect 33784 20757 33793 20791
rect 33793 20757 33827 20791
rect 33827 20757 33836 20791
rect 34152 20791 34204 20800
rect 33784 20748 33836 20757
rect 34152 20757 34161 20791
rect 34161 20757 34195 20791
rect 34195 20757 34204 20791
rect 34152 20748 34204 20757
rect 34980 20748 35032 20800
rect 4874 20646 4926 20698
rect 4938 20646 4990 20698
rect 5002 20646 5054 20698
rect 5066 20646 5118 20698
rect 5130 20646 5182 20698
rect 35594 20646 35646 20698
rect 35658 20646 35710 20698
rect 35722 20646 35774 20698
rect 35786 20646 35838 20698
rect 35850 20646 35902 20698
rect 7104 20544 7156 20596
rect 8668 20544 8720 20596
rect 11520 20544 11572 20596
rect 12900 20544 12952 20596
rect 13452 20587 13504 20596
rect 6828 20476 6880 20528
rect 8300 20476 8352 20528
rect 9956 20476 10008 20528
rect 11612 20476 11664 20528
rect 12440 20476 12492 20528
rect 13452 20553 13461 20587
rect 13461 20553 13495 20587
rect 13495 20553 13504 20587
rect 13452 20544 13504 20553
rect 15660 20544 15712 20596
rect 15936 20544 15988 20596
rect 17408 20544 17460 20596
rect 19432 20544 19484 20596
rect 25596 20587 25648 20596
rect 25596 20553 25605 20587
rect 25605 20553 25639 20587
rect 25639 20553 25648 20587
rect 25596 20544 25648 20553
rect 28172 20544 28224 20596
rect 29184 20544 29236 20596
rect 14464 20476 14516 20528
rect 15384 20476 15436 20528
rect 2136 20408 2188 20460
rect 8484 20451 8536 20460
rect 1584 20315 1636 20324
rect 1584 20281 1593 20315
rect 1593 20281 1627 20315
rect 1627 20281 1636 20315
rect 1584 20272 1636 20281
rect 8484 20417 8493 20451
rect 8493 20417 8527 20451
rect 8527 20417 8536 20451
rect 8484 20408 8536 20417
rect 9128 20408 9180 20460
rect 10784 20408 10836 20460
rect 11704 20451 11756 20460
rect 11704 20417 11713 20451
rect 11713 20417 11747 20451
rect 11747 20417 11756 20451
rect 11704 20408 11756 20417
rect 21824 20476 21876 20528
rect 24676 20476 24728 20528
rect 25320 20476 25372 20528
rect 30472 20544 30524 20596
rect 31576 20544 31628 20596
rect 35348 20544 35400 20596
rect 17776 20408 17828 20460
rect 10692 20340 10744 20392
rect 14096 20383 14148 20392
rect 14096 20349 14105 20383
rect 14105 20349 14139 20383
rect 14139 20349 14148 20383
rect 14096 20340 14148 20349
rect 20628 20451 20680 20460
rect 20628 20417 20637 20451
rect 20637 20417 20671 20451
rect 20671 20417 20680 20451
rect 20628 20408 20680 20417
rect 21180 20408 21232 20460
rect 22560 20451 22612 20460
rect 22560 20417 22569 20451
rect 22569 20417 22603 20451
rect 22603 20417 22612 20451
rect 22560 20408 22612 20417
rect 19800 20383 19852 20392
rect 19800 20349 19809 20383
rect 19809 20349 19843 20383
rect 19843 20349 19852 20383
rect 19800 20340 19852 20349
rect 20720 20340 20772 20392
rect 22008 20340 22060 20392
rect 24584 20340 24636 20392
rect 25780 20383 25832 20392
rect 25780 20349 25789 20383
rect 25789 20349 25823 20383
rect 25823 20349 25832 20383
rect 25780 20340 25832 20349
rect 27252 20340 27304 20392
rect 28724 20408 28776 20460
rect 30380 20408 30432 20460
rect 30840 20451 30892 20460
rect 30840 20417 30849 20451
rect 30849 20417 30883 20451
rect 30883 20417 30892 20451
rect 30840 20408 30892 20417
rect 31576 20408 31628 20460
rect 32864 20408 32916 20460
rect 34152 20408 34204 20460
rect 34980 20451 35032 20460
rect 34980 20417 34989 20451
rect 34989 20417 35023 20451
rect 35023 20417 35032 20451
rect 34980 20408 35032 20417
rect 36084 20476 36136 20528
rect 36636 20408 36688 20460
rect 29736 20383 29788 20392
rect 29736 20349 29745 20383
rect 29745 20349 29779 20383
rect 29779 20349 29788 20383
rect 33416 20383 33468 20392
rect 29736 20340 29788 20349
rect 33416 20349 33425 20383
rect 33425 20349 33459 20383
rect 33459 20349 33468 20383
rect 33416 20340 33468 20349
rect 33784 20340 33836 20392
rect 17592 20247 17644 20256
rect 17592 20213 17601 20247
rect 17601 20213 17635 20247
rect 17635 20213 17644 20247
rect 17592 20204 17644 20213
rect 19156 20204 19208 20256
rect 20720 20204 20772 20256
rect 21272 20204 21324 20256
rect 22376 20247 22428 20256
rect 22376 20213 22385 20247
rect 22385 20213 22419 20247
rect 22419 20213 22428 20247
rect 22376 20204 22428 20213
rect 25228 20247 25280 20256
rect 25228 20213 25237 20247
rect 25237 20213 25271 20247
rect 25271 20213 25280 20247
rect 25228 20204 25280 20213
rect 26976 20204 27028 20256
rect 30564 20272 30616 20324
rect 36912 20315 36964 20324
rect 36912 20281 36921 20315
rect 36921 20281 36955 20315
rect 36955 20281 36964 20315
rect 36912 20272 36964 20281
rect 28264 20204 28316 20256
rect 31300 20247 31352 20256
rect 31300 20213 31309 20247
rect 31309 20213 31343 20247
rect 31343 20213 31352 20247
rect 31300 20204 31352 20213
rect 34060 20204 34112 20256
rect 35716 20247 35768 20256
rect 35716 20213 35725 20247
rect 35725 20213 35759 20247
rect 35759 20213 35768 20247
rect 35716 20204 35768 20213
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 10140 20000 10192 20052
rect 12440 20043 12492 20052
rect 12440 20009 12449 20043
rect 12449 20009 12483 20043
rect 12483 20009 12492 20043
rect 14280 20043 14332 20052
rect 12440 20000 12492 20009
rect 14280 20009 14289 20043
rect 14289 20009 14323 20043
rect 14323 20009 14332 20043
rect 14280 20000 14332 20009
rect 19708 20000 19760 20052
rect 14740 19932 14792 19984
rect 16028 19932 16080 19984
rect 17684 19932 17736 19984
rect 11060 19864 11112 19916
rect 11520 19907 11572 19916
rect 11520 19873 11529 19907
rect 11529 19873 11563 19907
rect 11563 19873 11572 19907
rect 11520 19864 11572 19873
rect 12808 19864 12860 19916
rect 13084 19907 13136 19916
rect 13084 19873 13093 19907
rect 13093 19873 13127 19907
rect 13127 19873 13136 19907
rect 13084 19864 13136 19873
rect 8576 19839 8628 19848
rect 8576 19805 8585 19839
rect 8585 19805 8619 19839
rect 8619 19805 8628 19839
rect 8576 19796 8628 19805
rect 9496 19796 9548 19848
rect 12164 19796 12216 19848
rect 12440 19796 12492 19848
rect 13452 19796 13504 19848
rect 15936 19864 15988 19916
rect 21180 20000 21232 20052
rect 22284 20000 22336 20052
rect 22560 20000 22612 20052
rect 24584 20043 24636 20052
rect 24584 20009 24593 20043
rect 24593 20009 24627 20043
rect 24627 20009 24636 20043
rect 24584 20000 24636 20009
rect 28172 20000 28224 20052
rect 32496 20000 32548 20052
rect 15660 19839 15712 19848
rect 15660 19805 15669 19839
rect 15669 19805 15703 19839
rect 15703 19805 15712 19839
rect 15660 19796 15712 19805
rect 18696 19839 18748 19848
rect 18696 19805 18705 19839
rect 18705 19805 18739 19839
rect 18739 19805 18748 19839
rect 22008 19864 22060 19916
rect 25136 19932 25188 19984
rect 18696 19796 18748 19805
rect 18880 19796 18932 19848
rect 25228 19864 25280 19916
rect 25320 19864 25372 19916
rect 26976 19907 27028 19916
rect 26976 19873 26985 19907
rect 26985 19873 27019 19907
rect 27019 19873 27028 19907
rect 26976 19864 27028 19873
rect 31208 19864 31260 19916
rect 34060 19907 34112 19916
rect 34060 19873 34069 19907
rect 34069 19873 34103 19907
rect 34103 19873 34112 19907
rect 34060 19864 34112 19873
rect 34336 19907 34388 19916
rect 34336 19873 34345 19907
rect 34345 19873 34379 19907
rect 34379 19873 34388 19907
rect 34336 19864 34388 19873
rect 24768 19839 24820 19848
rect 24768 19805 24777 19839
rect 24777 19805 24811 19839
rect 24811 19805 24820 19839
rect 24768 19796 24820 19805
rect 26424 19796 26476 19848
rect 9588 19728 9640 19780
rect 11612 19728 11664 19780
rect 14464 19728 14516 19780
rect 8392 19703 8444 19712
rect 8392 19669 8401 19703
rect 8401 19669 8435 19703
rect 8435 19669 8444 19703
rect 8392 19660 8444 19669
rect 9312 19660 9364 19712
rect 10600 19660 10652 19712
rect 13728 19703 13780 19712
rect 13728 19669 13737 19703
rect 13737 19669 13771 19703
rect 13771 19669 13780 19703
rect 13728 19660 13780 19669
rect 17592 19728 17644 19780
rect 20720 19771 20772 19780
rect 20720 19737 20729 19771
rect 20729 19737 20763 19771
rect 20763 19737 20772 19771
rect 20720 19728 20772 19737
rect 21272 19728 21324 19780
rect 17960 19660 18012 19712
rect 18788 19703 18840 19712
rect 18788 19669 18797 19703
rect 18797 19669 18831 19703
rect 18831 19669 18840 19703
rect 18788 19660 18840 19669
rect 18972 19660 19024 19712
rect 23756 19703 23808 19712
rect 23756 19669 23765 19703
rect 23765 19669 23799 19703
rect 23799 19669 23808 19703
rect 23756 19660 23808 19669
rect 25044 19660 25096 19712
rect 25872 19703 25924 19712
rect 25872 19669 25881 19703
rect 25881 19669 25915 19703
rect 25915 19669 25924 19703
rect 25872 19660 25924 19669
rect 26792 19660 26844 19712
rect 28264 19728 28316 19780
rect 30840 19728 30892 19780
rect 31300 19771 31352 19780
rect 31300 19737 31309 19771
rect 31309 19737 31343 19771
rect 31343 19737 31352 19771
rect 31300 19728 31352 19737
rect 35716 19728 35768 19780
rect 29736 19660 29788 19712
rect 4874 19558 4926 19610
rect 4938 19558 4990 19610
rect 5002 19558 5054 19610
rect 5066 19558 5118 19610
rect 5130 19558 5182 19610
rect 35594 19558 35646 19610
rect 35658 19558 35710 19610
rect 35722 19558 35774 19610
rect 35786 19558 35838 19610
rect 35850 19558 35902 19610
rect 8576 19456 8628 19508
rect 10600 19499 10652 19508
rect 10600 19465 10609 19499
rect 10609 19465 10643 19499
rect 10643 19465 10652 19499
rect 10600 19456 10652 19465
rect 8300 19388 8352 19440
rect 9312 19388 9364 19440
rect 9588 19320 9640 19372
rect 8392 19252 8444 19304
rect 11888 19363 11940 19372
rect 11888 19329 11897 19363
rect 11897 19329 11931 19363
rect 11931 19329 11940 19363
rect 11888 19320 11940 19329
rect 13728 19456 13780 19508
rect 15660 19456 15712 19508
rect 18972 19456 19024 19508
rect 20628 19499 20680 19508
rect 20628 19465 20637 19499
rect 20637 19465 20671 19499
rect 20671 19465 20680 19499
rect 20628 19456 20680 19465
rect 20812 19456 20864 19508
rect 22284 19456 22336 19508
rect 23756 19456 23808 19508
rect 12624 19388 12676 19440
rect 14096 19388 14148 19440
rect 14464 19320 14516 19372
rect 15292 19388 15344 19440
rect 18880 19388 18932 19440
rect 21088 19431 21140 19440
rect 21088 19397 21097 19431
rect 21097 19397 21131 19431
rect 21131 19397 21140 19431
rect 21088 19388 21140 19397
rect 22376 19431 22428 19440
rect 22376 19397 22385 19431
rect 22385 19397 22419 19431
rect 22419 19397 22428 19431
rect 22376 19388 22428 19397
rect 24308 19388 24360 19440
rect 19892 19363 19944 19372
rect 19892 19329 19901 19363
rect 19901 19329 19935 19363
rect 19935 19329 19944 19363
rect 19892 19320 19944 19329
rect 22008 19320 22060 19372
rect 25044 19431 25096 19440
rect 25044 19397 25053 19431
rect 25053 19397 25087 19431
rect 25087 19397 25096 19431
rect 25044 19388 25096 19397
rect 27252 19456 27304 19508
rect 29000 19456 29052 19508
rect 30840 19499 30892 19508
rect 30840 19465 30849 19499
rect 30849 19465 30883 19499
rect 30883 19465 30892 19499
rect 30840 19456 30892 19465
rect 10692 19184 10744 19236
rect 12716 19252 12768 19304
rect 13636 19252 13688 19304
rect 13728 19252 13780 19304
rect 17316 19295 17368 19304
rect 17316 19261 17325 19295
rect 17325 19261 17359 19295
rect 17359 19261 17368 19295
rect 17316 19252 17368 19261
rect 16488 19184 16540 19236
rect 19156 19252 19208 19304
rect 20260 19252 20312 19304
rect 25136 19295 25188 19304
rect 25136 19261 25145 19295
rect 25145 19261 25179 19295
rect 25179 19261 25188 19295
rect 25136 19252 25188 19261
rect 25872 19252 25924 19304
rect 32772 19388 32824 19440
rect 26424 19320 26476 19372
rect 28724 19320 28776 19372
rect 30564 19320 30616 19372
rect 31576 19320 31628 19372
rect 34336 19320 34388 19372
rect 25780 19184 25832 19236
rect 26976 19252 27028 19304
rect 31024 19252 31076 19304
rect 11704 19159 11756 19168
rect 11704 19125 11713 19159
rect 11713 19125 11747 19159
rect 11747 19125 11756 19159
rect 11704 19116 11756 19125
rect 12900 19116 12952 19168
rect 18052 19116 18104 19168
rect 23940 19116 23992 19168
rect 28448 19116 28500 19168
rect 31392 19116 31444 19168
rect 31852 19116 31904 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 1768 18912 1820 18964
rect 7012 18912 7064 18964
rect 11888 18912 11940 18964
rect 13728 18955 13780 18964
rect 13728 18921 13737 18955
rect 13737 18921 13771 18955
rect 13771 18921 13780 18955
rect 13728 18912 13780 18921
rect 15292 18912 15344 18964
rect 15660 18912 15712 18964
rect 18880 18912 18932 18964
rect 19432 18955 19484 18964
rect 19432 18921 19441 18955
rect 19441 18921 19475 18955
rect 19475 18921 19484 18955
rect 19432 18912 19484 18921
rect 25044 18912 25096 18964
rect 26976 18955 27028 18964
rect 26976 18921 26985 18955
rect 26985 18921 27019 18955
rect 27019 18921 27028 18955
rect 26976 18912 27028 18921
rect 31024 18955 31076 18964
rect 31024 18921 31033 18955
rect 31033 18921 31067 18955
rect 31067 18921 31076 18955
rect 31024 18912 31076 18921
rect 32772 18912 32824 18964
rect 16580 18844 16632 18896
rect 19800 18844 19852 18896
rect 8300 18776 8352 18828
rect 9404 18776 9456 18828
rect 11060 18776 11112 18828
rect 11612 18819 11664 18828
rect 11612 18785 11621 18819
rect 11621 18785 11655 18819
rect 11655 18785 11664 18819
rect 11612 18776 11664 18785
rect 12440 18776 12492 18828
rect 13728 18776 13780 18828
rect 16212 18776 16264 18828
rect 16948 18776 17000 18828
rect 6000 18640 6052 18692
rect 7288 18640 7340 18692
rect 8392 18640 8444 18692
rect 9864 18640 9916 18692
rect 13544 18751 13596 18760
rect 13544 18717 13553 18751
rect 13553 18717 13587 18751
rect 13587 18717 13596 18751
rect 13544 18708 13596 18717
rect 14280 18751 14332 18760
rect 14280 18717 14289 18751
rect 14289 18717 14323 18751
rect 14323 18717 14332 18751
rect 14280 18708 14332 18717
rect 14464 18708 14516 18760
rect 16488 18751 16540 18760
rect 16488 18717 16497 18751
rect 16497 18717 16531 18751
rect 16531 18717 16540 18751
rect 16488 18708 16540 18717
rect 17316 18708 17368 18760
rect 13360 18640 13412 18692
rect 15476 18640 15528 18692
rect 20260 18776 20312 18828
rect 22008 18776 22060 18828
rect 30748 18819 30800 18828
rect 17776 18708 17828 18760
rect 22100 18751 22152 18760
rect 22100 18717 22109 18751
rect 22109 18717 22143 18751
rect 22143 18717 22152 18751
rect 22100 18708 22152 18717
rect 18788 18640 18840 18692
rect 20904 18683 20956 18692
rect 20904 18649 20913 18683
rect 20913 18649 20947 18683
rect 20947 18649 20956 18683
rect 20904 18640 20956 18649
rect 21916 18640 21968 18692
rect 23940 18708 23992 18760
rect 26792 18751 26844 18760
rect 26792 18717 26801 18751
rect 26801 18717 26835 18751
rect 26835 18717 26844 18751
rect 26792 18708 26844 18717
rect 27528 18708 27580 18760
rect 29000 18751 29052 18760
rect 29000 18717 29009 18751
rect 29009 18717 29043 18751
rect 29043 18717 29052 18751
rect 29000 18708 29052 18717
rect 29184 18751 29236 18760
rect 29184 18717 29193 18751
rect 29193 18717 29227 18751
rect 29227 18717 29236 18751
rect 29184 18708 29236 18717
rect 30748 18785 30757 18819
rect 30757 18785 30791 18819
rect 30791 18785 30800 18819
rect 30748 18776 30800 18785
rect 2044 18572 2096 18624
rect 9680 18572 9732 18624
rect 12164 18572 12216 18624
rect 12992 18615 13044 18624
rect 12992 18581 13001 18615
rect 13001 18581 13035 18615
rect 13035 18581 13044 18615
rect 12992 18572 13044 18581
rect 14924 18615 14976 18624
rect 14924 18581 14933 18615
rect 14933 18581 14967 18615
rect 14967 18581 14976 18615
rect 14924 18572 14976 18581
rect 15200 18572 15252 18624
rect 16580 18572 16632 18624
rect 17500 18615 17552 18624
rect 17500 18581 17509 18615
rect 17509 18581 17543 18615
rect 17543 18581 17552 18615
rect 22928 18615 22980 18624
rect 17500 18572 17552 18581
rect 22928 18581 22937 18615
rect 22937 18581 22971 18615
rect 22971 18581 22980 18615
rect 22928 18572 22980 18581
rect 25320 18640 25372 18692
rect 28356 18683 28408 18692
rect 28356 18649 28365 18683
rect 28365 18649 28399 18683
rect 28399 18649 28408 18683
rect 28356 18640 28408 18649
rect 31852 18708 31904 18760
rect 32312 18751 32364 18760
rect 32312 18717 32321 18751
rect 32321 18717 32355 18751
rect 32355 18717 32364 18751
rect 32312 18708 32364 18717
rect 33416 18708 33468 18760
rect 31300 18640 31352 18692
rect 28816 18572 28868 18624
rect 30288 18572 30340 18624
rect 35072 18572 35124 18624
rect 4874 18470 4926 18522
rect 4938 18470 4990 18522
rect 5002 18470 5054 18522
rect 5066 18470 5118 18522
rect 5130 18470 5182 18522
rect 35594 18470 35646 18522
rect 35658 18470 35710 18522
rect 35722 18470 35774 18522
rect 35786 18470 35838 18522
rect 35850 18470 35902 18522
rect 6000 18411 6052 18420
rect 6000 18377 6009 18411
rect 6009 18377 6043 18411
rect 6043 18377 6052 18411
rect 6000 18368 6052 18377
rect 7288 18368 7340 18420
rect 9864 18368 9916 18420
rect 11152 18411 11204 18420
rect 6368 18232 6420 18284
rect 7288 18275 7340 18284
rect 7288 18241 7297 18275
rect 7297 18241 7331 18275
rect 7331 18241 7340 18275
rect 9772 18300 9824 18352
rect 10140 18300 10192 18352
rect 11152 18377 11161 18411
rect 11161 18377 11195 18411
rect 11195 18377 11204 18411
rect 11152 18368 11204 18377
rect 11612 18368 11664 18420
rect 13544 18368 13596 18420
rect 15200 18411 15252 18420
rect 15200 18377 15209 18411
rect 15209 18377 15243 18411
rect 15243 18377 15252 18411
rect 15200 18368 15252 18377
rect 12900 18343 12952 18352
rect 7288 18232 7340 18241
rect 9220 18232 9272 18284
rect 9404 18275 9456 18284
rect 9404 18241 9413 18275
rect 9413 18241 9447 18275
rect 9447 18241 9456 18275
rect 9404 18232 9456 18241
rect 12900 18309 12909 18343
rect 12909 18309 12943 18343
rect 12943 18309 12952 18343
rect 12900 18300 12952 18309
rect 12992 18300 13044 18352
rect 19432 18411 19484 18420
rect 19432 18377 19441 18411
rect 19441 18377 19475 18411
rect 19475 18377 19484 18411
rect 19432 18368 19484 18377
rect 20812 18411 20864 18420
rect 20812 18377 20821 18411
rect 20821 18377 20855 18411
rect 20855 18377 20864 18411
rect 20812 18368 20864 18377
rect 21916 18368 21968 18420
rect 16580 18300 16632 18352
rect 18144 18300 18196 18352
rect 12624 18207 12676 18216
rect 12624 18173 12633 18207
rect 12633 18173 12667 18207
rect 12667 18173 12676 18207
rect 12624 18164 12676 18173
rect 14464 18164 14516 18216
rect 15292 18207 15344 18216
rect 15292 18173 15301 18207
rect 15301 18173 15335 18207
rect 15335 18173 15344 18207
rect 15292 18164 15344 18173
rect 15476 18207 15528 18216
rect 15476 18173 15485 18207
rect 15485 18173 15519 18207
rect 15519 18173 15528 18207
rect 15476 18164 15528 18173
rect 16764 18164 16816 18216
rect 20904 18300 20956 18352
rect 22928 18300 22980 18352
rect 20720 18275 20772 18284
rect 20720 18241 20729 18275
rect 20729 18241 20763 18275
rect 20763 18241 20772 18275
rect 20720 18232 20772 18241
rect 25320 18368 25372 18420
rect 25044 18300 25096 18352
rect 26056 18275 26108 18284
rect 26056 18241 26065 18275
rect 26065 18241 26099 18275
rect 26099 18241 26108 18275
rect 26056 18232 26108 18241
rect 26792 18232 26844 18284
rect 29460 18368 29512 18420
rect 20260 18164 20312 18216
rect 20996 18207 21048 18216
rect 20996 18173 21005 18207
rect 21005 18173 21039 18207
rect 21039 18173 21048 18207
rect 20996 18164 21048 18173
rect 22008 18207 22060 18216
rect 22008 18173 22017 18207
rect 22017 18173 22051 18207
rect 22051 18173 22060 18207
rect 22008 18164 22060 18173
rect 22284 18207 22336 18216
rect 22284 18173 22293 18207
rect 22293 18173 22327 18207
rect 22327 18173 22336 18207
rect 22284 18164 22336 18173
rect 25320 18207 25372 18216
rect 25320 18173 25329 18207
rect 25329 18173 25363 18207
rect 25363 18173 25372 18207
rect 25320 18164 25372 18173
rect 25504 18207 25556 18216
rect 25504 18173 25513 18207
rect 25513 18173 25547 18207
rect 25547 18173 25556 18207
rect 25504 18164 25556 18173
rect 25780 18164 25832 18216
rect 26976 18164 27028 18216
rect 27528 18300 27580 18352
rect 28816 18343 28868 18352
rect 28816 18309 28825 18343
rect 28825 18309 28859 18343
rect 28859 18309 28868 18343
rect 28816 18300 28868 18309
rect 31208 18368 31260 18420
rect 31760 18411 31812 18420
rect 31760 18377 31769 18411
rect 31769 18377 31803 18411
rect 31803 18377 31812 18411
rect 31760 18368 31812 18377
rect 30288 18343 30340 18352
rect 28540 18275 28592 18284
rect 28540 18241 28549 18275
rect 28549 18241 28583 18275
rect 28583 18241 28592 18275
rect 28540 18232 28592 18241
rect 28632 18275 28684 18284
rect 28632 18241 28642 18275
rect 28642 18241 28676 18275
rect 28676 18241 28684 18275
rect 28632 18232 28684 18241
rect 28080 18164 28132 18216
rect 29092 18232 29144 18284
rect 30288 18309 30297 18343
rect 30297 18309 30331 18343
rect 30331 18309 30340 18343
rect 30288 18300 30340 18309
rect 32404 18368 32456 18420
rect 30380 18164 30432 18216
rect 33416 18232 33468 18284
rect 34336 18300 34388 18352
rect 35072 18300 35124 18352
rect 34060 18207 34112 18216
rect 34060 18173 34069 18207
rect 34069 18173 34103 18207
rect 34103 18173 34112 18207
rect 34060 18164 34112 18173
rect 31300 18096 31352 18148
rect 12072 18071 12124 18080
rect 12072 18037 12081 18071
rect 12081 18037 12115 18071
rect 12115 18037 12124 18071
rect 12072 18028 12124 18037
rect 17316 18028 17368 18080
rect 20352 18071 20404 18080
rect 20352 18037 20361 18071
rect 20361 18037 20395 18071
rect 20395 18037 20404 18071
rect 20352 18028 20404 18037
rect 23664 18028 23716 18080
rect 24860 18071 24912 18080
rect 24860 18037 24869 18071
rect 24869 18037 24903 18071
rect 24903 18037 24912 18071
rect 24860 18028 24912 18037
rect 26700 18028 26752 18080
rect 29460 18028 29512 18080
rect 30932 18028 30984 18080
rect 31760 18028 31812 18080
rect 34796 18028 34848 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 8392 17824 8444 17876
rect 10140 17824 10192 17876
rect 12164 17824 12216 17876
rect 18052 17824 18104 17876
rect 22284 17824 22336 17876
rect 26056 17824 26108 17876
rect 28632 17867 28684 17876
rect 28632 17833 28641 17867
rect 28641 17833 28675 17867
rect 28675 17833 28684 17867
rect 28632 17824 28684 17833
rect 34060 17824 34112 17876
rect 13360 17756 13412 17808
rect 16028 17799 16080 17808
rect 16028 17765 16037 17799
rect 16037 17765 16071 17799
rect 16071 17765 16080 17799
rect 16028 17756 16080 17765
rect 7104 17731 7156 17740
rect 7104 17697 7113 17731
rect 7113 17697 7147 17731
rect 7147 17697 7156 17731
rect 7104 17688 7156 17697
rect 10692 17731 10744 17740
rect 10692 17697 10701 17731
rect 10701 17697 10735 17731
rect 10735 17697 10744 17731
rect 10692 17688 10744 17697
rect 12624 17688 12676 17740
rect 13636 17688 13688 17740
rect 15292 17688 15344 17740
rect 16948 17731 17000 17740
rect 16948 17697 16957 17731
rect 16957 17697 16991 17731
rect 16991 17697 17000 17731
rect 16948 17688 17000 17697
rect 17316 17688 17368 17740
rect 19432 17688 19484 17740
rect 6092 17552 6144 17604
rect 6644 17552 6696 17604
rect 8760 17620 8812 17672
rect 9496 17663 9548 17672
rect 9496 17629 9505 17663
rect 9505 17629 9539 17663
rect 9539 17629 9548 17663
rect 9496 17620 9548 17629
rect 11152 17620 11204 17672
rect 14924 17620 14976 17672
rect 18696 17620 18748 17672
rect 20352 17663 20404 17672
rect 20352 17629 20361 17663
rect 20361 17629 20395 17663
rect 20395 17629 20404 17663
rect 20352 17620 20404 17629
rect 23664 17731 23716 17740
rect 23664 17697 23673 17731
rect 23673 17697 23707 17731
rect 23707 17697 23716 17731
rect 23664 17688 23716 17697
rect 21916 17663 21968 17672
rect 21916 17629 21925 17663
rect 21925 17629 21959 17663
rect 21959 17629 21968 17663
rect 21916 17620 21968 17629
rect 10784 17552 10836 17604
rect 11704 17552 11756 17604
rect 12072 17552 12124 17604
rect 16304 17595 16356 17604
rect 16304 17561 16313 17595
rect 16313 17561 16347 17595
rect 16347 17561 16356 17595
rect 16304 17552 16356 17561
rect 17132 17552 17184 17604
rect 17500 17552 17552 17604
rect 18604 17552 18656 17604
rect 21088 17552 21140 17604
rect 6736 17484 6788 17536
rect 6920 17527 6972 17536
rect 6920 17493 6929 17527
rect 6929 17493 6963 17527
rect 6963 17493 6972 17527
rect 6920 17484 6972 17493
rect 9220 17484 9272 17536
rect 10508 17527 10560 17536
rect 10508 17493 10517 17527
rect 10517 17493 10551 17527
rect 10551 17493 10560 17527
rect 10508 17484 10560 17493
rect 15384 17484 15436 17536
rect 16488 17484 16540 17536
rect 17592 17527 17644 17536
rect 17592 17493 17601 17527
rect 17601 17493 17635 17527
rect 17635 17493 17644 17527
rect 17592 17484 17644 17493
rect 18880 17527 18932 17536
rect 18880 17493 18889 17527
rect 18889 17493 18923 17527
rect 18923 17493 18932 17527
rect 18880 17484 18932 17493
rect 21180 17527 21232 17536
rect 21180 17493 21189 17527
rect 21189 17493 21223 17527
rect 21223 17493 21232 17527
rect 21180 17484 21232 17493
rect 22744 17484 22796 17536
rect 23388 17620 23440 17672
rect 25136 17688 25188 17740
rect 25228 17688 25280 17740
rect 26700 17731 26752 17740
rect 26700 17697 26709 17731
rect 26709 17697 26743 17731
rect 26743 17697 26752 17731
rect 26700 17688 26752 17697
rect 30380 17688 30432 17740
rect 31208 17731 31260 17740
rect 31208 17697 31217 17731
rect 31217 17697 31251 17731
rect 31251 17697 31260 17731
rect 31208 17688 31260 17697
rect 32680 17688 32732 17740
rect 34796 17688 34848 17740
rect 25412 17620 25464 17672
rect 26424 17663 26476 17672
rect 26424 17629 26433 17663
rect 26433 17629 26467 17663
rect 26467 17629 26476 17663
rect 26424 17620 26476 17629
rect 27804 17620 27856 17672
rect 28908 17620 28960 17672
rect 29184 17620 29236 17672
rect 29920 17663 29972 17672
rect 29920 17629 29929 17663
rect 29929 17629 29963 17663
rect 29963 17629 29972 17663
rect 29920 17620 29972 17629
rect 32956 17663 33008 17672
rect 32956 17629 32965 17663
rect 32965 17629 32999 17663
rect 32999 17629 33008 17663
rect 32956 17620 33008 17629
rect 34060 17620 34112 17672
rect 24860 17552 24912 17604
rect 25320 17552 25372 17604
rect 24768 17527 24820 17536
rect 24768 17493 24777 17527
rect 24777 17493 24811 17527
rect 24811 17493 24820 17527
rect 24768 17484 24820 17493
rect 35072 17552 35124 17604
rect 35348 17552 35400 17604
rect 28172 17527 28224 17536
rect 28172 17493 28181 17527
rect 28181 17493 28215 17527
rect 28215 17493 28224 17527
rect 28172 17484 28224 17493
rect 30288 17527 30340 17536
rect 30288 17493 30297 17527
rect 30297 17493 30331 17527
rect 30331 17493 30340 17527
rect 30288 17484 30340 17493
rect 35256 17484 35308 17536
rect 4874 17382 4926 17434
rect 4938 17382 4990 17434
rect 5002 17382 5054 17434
rect 5066 17382 5118 17434
rect 5130 17382 5182 17434
rect 35594 17382 35646 17434
rect 35658 17382 35710 17434
rect 35722 17382 35774 17434
rect 35786 17382 35838 17434
rect 35850 17382 35902 17434
rect 8208 17280 8260 17332
rect 8760 17323 8812 17332
rect 8760 17289 8769 17323
rect 8769 17289 8803 17323
rect 8803 17289 8812 17323
rect 8760 17280 8812 17289
rect 9680 17280 9732 17332
rect 10508 17280 10560 17332
rect 12164 17323 12216 17332
rect 12164 17289 12173 17323
rect 12173 17289 12207 17323
rect 12207 17289 12216 17323
rect 12164 17280 12216 17289
rect 13636 17280 13688 17332
rect 5816 17187 5868 17196
rect 5816 17153 5825 17187
rect 5825 17153 5859 17187
rect 5859 17153 5868 17187
rect 5816 17144 5868 17153
rect 6092 17144 6144 17196
rect 6552 17119 6604 17128
rect 6552 17085 6561 17119
rect 6561 17085 6595 17119
rect 6595 17085 6604 17119
rect 6552 17076 6604 17085
rect 6828 17119 6880 17128
rect 6828 17085 6837 17119
rect 6837 17085 6871 17119
rect 6871 17085 6880 17119
rect 6828 17076 6880 17085
rect 1584 16983 1636 16992
rect 1584 16949 1593 16983
rect 1593 16949 1627 16983
rect 1627 16949 1636 16983
rect 1584 16940 1636 16949
rect 6828 16940 6880 16992
rect 15568 17212 15620 17264
rect 12440 17144 12492 17196
rect 14096 17144 14148 17196
rect 9220 17119 9272 17128
rect 9220 17085 9229 17119
rect 9229 17085 9263 17119
rect 9263 17085 9272 17119
rect 9220 17076 9272 17085
rect 10600 17119 10652 17128
rect 9036 17008 9088 17060
rect 10600 17085 10609 17119
rect 10609 17085 10643 17119
rect 10643 17085 10652 17119
rect 10600 17076 10652 17085
rect 12900 17076 12952 17128
rect 13360 17076 13412 17128
rect 14832 17119 14884 17128
rect 13268 17008 13320 17060
rect 14832 17085 14841 17119
rect 14841 17085 14875 17119
rect 14875 17085 14884 17119
rect 14832 17076 14884 17085
rect 15292 17076 15344 17128
rect 16488 17076 16540 17128
rect 17592 17280 17644 17332
rect 18880 17323 18932 17332
rect 18880 17289 18889 17323
rect 18889 17289 18923 17323
rect 18923 17289 18932 17323
rect 18880 17280 18932 17289
rect 21088 17280 21140 17332
rect 23664 17280 23716 17332
rect 25412 17323 25464 17332
rect 25412 17289 25421 17323
rect 25421 17289 25455 17323
rect 25455 17289 25464 17323
rect 25412 17280 25464 17289
rect 28540 17280 28592 17332
rect 17500 17212 17552 17264
rect 20444 17212 20496 17264
rect 21180 17255 21232 17264
rect 21180 17221 21189 17255
rect 21189 17221 21223 17255
rect 21223 17221 21232 17255
rect 21180 17212 21232 17221
rect 22744 17212 22796 17264
rect 29920 17280 29972 17332
rect 30380 17280 30432 17332
rect 31208 17280 31260 17332
rect 30288 17255 30340 17264
rect 27252 17144 27304 17196
rect 18696 17076 18748 17128
rect 20720 17076 20772 17128
rect 21640 17076 21692 17128
rect 22008 17119 22060 17128
rect 22008 17085 22017 17119
rect 22017 17085 22051 17119
rect 22051 17085 22060 17119
rect 22008 17076 22060 17085
rect 22284 17119 22336 17128
rect 22284 17085 22293 17119
rect 22293 17085 22327 17119
rect 22327 17085 22336 17119
rect 22284 17076 22336 17085
rect 24952 17076 25004 17128
rect 25504 17076 25556 17128
rect 9956 16983 10008 16992
rect 9956 16949 9965 16983
rect 9965 16949 9999 16983
rect 9999 16949 10008 16983
rect 9956 16940 10008 16949
rect 13636 16983 13688 16992
rect 13636 16949 13645 16983
rect 13645 16949 13679 16983
rect 13679 16949 13688 16983
rect 13636 16940 13688 16949
rect 16764 17008 16816 17060
rect 23480 17008 23532 17060
rect 24584 17008 24636 17060
rect 16948 16940 17000 16992
rect 18880 16940 18932 16992
rect 24216 16983 24268 16992
rect 24216 16949 24225 16983
rect 24225 16949 24259 16983
rect 24259 16949 24268 16983
rect 24216 16940 24268 16949
rect 25228 16940 25280 16992
rect 25504 16940 25556 16992
rect 27160 17076 27212 17128
rect 29000 17144 29052 17196
rect 30288 17221 30297 17255
rect 30297 17221 30331 17255
rect 30331 17221 30340 17255
rect 30288 17212 30340 17221
rect 31668 17212 31720 17264
rect 34336 17280 34388 17332
rect 35072 17280 35124 17332
rect 35440 17280 35492 17332
rect 33232 17212 33284 17264
rect 35256 17212 35308 17264
rect 35900 17212 35952 17264
rect 28080 17076 28132 17128
rect 27068 16940 27120 16992
rect 34336 17144 34388 17196
rect 33324 17076 33376 17128
rect 34060 17119 34112 17128
rect 34060 17085 34069 17119
rect 34069 17085 34103 17119
rect 34103 17085 34112 17119
rect 34060 17076 34112 17085
rect 31852 16940 31904 16992
rect 32404 16940 32456 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 7104 16736 7156 16788
rect 9588 16736 9640 16788
rect 10692 16736 10744 16788
rect 13728 16736 13780 16788
rect 18604 16779 18656 16788
rect 18604 16745 18613 16779
rect 18613 16745 18647 16779
rect 18647 16745 18656 16779
rect 18604 16736 18656 16745
rect 20720 16736 20772 16788
rect 22284 16779 22336 16788
rect 22284 16745 22293 16779
rect 22293 16745 22327 16779
rect 22327 16745 22336 16779
rect 22284 16736 22336 16745
rect 24768 16736 24820 16788
rect 27252 16779 27304 16788
rect 27252 16745 27261 16779
rect 27261 16745 27295 16779
rect 27295 16745 27304 16779
rect 27252 16736 27304 16745
rect 27620 16736 27672 16788
rect 29184 16736 29236 16788
rect 30748 16779 30800 16788
rect 30748 16745 30757 16779
rect 30757 16745 30791 16779
rect 30791 16745 30800 16779
rect 30748 16736 30800 16745
rect 30932 16779 30984 16788
rect 30932 16745 30941 16779
rect 30941 16745 30975 16779
rect 30975 16745 30984 16779
rect 30932 16736 30984 16745
rect 34796 16736 34848 16788
rect 35348 16736 35400 16788
rect 35900 16736 35952 16788
rect 6092 16668 6144 16720
rect 6828 16643 6880 16652
rect 6828 16609 6837 16643
rect 6837 16609 6871 16643
rect 6871 16609 6880 16643
rect 6828 16600 6880 16609
rect 7196 16600 7248 16652
rect 8208 16643 8260 16652
rect 7012 16532 7064 16584
rect 8208 16609 8217 16643
rect 8217 16609 8251 16643
rect 8251 16609 8260 16643
rect 8208 16600 8260 16609
rect 14096 16668 14148 16720
rect 23388 16668 23440 16720
rect 24952 16711 25004 16720
rect 12900 16643 12952 16652
rect 12900 16609 12909 16643
rect 12909 16609 12943 16643
rect 12943 16609 12952 16643
rect 12900 16600 12952 16609
rect 13360 16600 13412 16652
rect 14280 16600 14332 16652
rect 10784 16532 10836 16584
rect 13636 16575 13688 16584
rect 6644 16464 6696 16516
rect 9404 16507 9456 16516
rect 6368 16439 6420 16448
rect 6368 16405 6377 16439
rect 6377 16405 6411 16439
rect 6411 16405 6420 16439
rect 6368 16396 6420 16405
rect 9404 16473 9413 16507
rect 9413 16473 9447 16507
rect 9447 16473 9456 16507
rect 9404 16464 9456 16473
rect 10140 16464 10192 16516
rect 7932 16439 7984 16448
rect 7932 16405 7941 16439
rect 7941 16405 7975 16439
rect 7975 16405 7984 16439
rect 7932 16396 7984 16405
rect 9220 16396 9272 16448
rect 13636 16541 13645 16575
rect 13645 16541 13679 16575
rect 13679 16541 13688 16575
rect 13636 16532 13688 16541
rect 14648 16575 14700 16584
rect 14648 16541 14657 16575
rect 14657 16541 14691 16575
rect 14691 16541 14700 16575
rect 14648 16532 14700 16541
rect 15660 16532 15712 16584
rect 16764 16600 16816 16652
rect 21640 16600 21692 16652
rect 23480 16643 23532 16652
rect 23480 16609 23489 16643
rect 23489 16609 23523 16643
rect 23523 16609 23532 16643
rect 23480 16600 23532 16609
rect 24952 16677 24961 16711
rect 24961 16677 24995 16711
rect 24995 16677 25004 16711
rect 24952 16668 25004 16677
rect 26424 16600 26476 16652
rect 27160 16600 27212 16652
rect 28724 16668 28776 16720
rect 29000 16668 29052 16720
rect 14464 16464 14516 16516
rect 11980 16396 12032 16448
rect 12256 16439 12308 16448
rect 12256 16405 12265 16439
rect 12265 16405 12299 16439
rect 12299 16405 12308 16439
rect 12256 16396 12308 16405
rect 13544 16396 13596 16448
rect 16580 16464 16632 16516
rect 17132 16507 17184 16516
rect 17132 16473 17141 16507
rect 17141 16473 17175 16507
rect 17175 16473 17184 16507
rect 17132 16464 17184 16473
rect 18144 16464 18196 16516
rect 19340 16464 19392 16516
rect 20168 16464 20220 16516
rect 18052 16396 18104 16448
rect 24216 16532 24268 16584
rect 27804 16575 27856 16584
rect 27804 16541 27813 16575
rect 27813 16541 27847 16575
rect 27847 16541 27856 16575
rect 27804 16532 27856 16541
rect 28172 16600 28224 16652
rect 29736 16575 29788 16584
rect 29736 16541 29745 16575
rect 29745 16541 29779 16575
rect 29779 16541 29788 16575
rect 29736 16532 29788 16541
rect 30012 16575 30064 16584
rect 30012 16541 30021 16575
rect 30021 16541 30055 16575
rect 30055 16541 30064 16575
rect 30012 16532 30064 16541
rect 31668 16575 31720 16584
rect 31668 16541 31677 16575
rect 31677 16541 31711 16575
rect 31711 16541 31720 16575
rect 31668 16532 31720 16541
rect 32680 16575 32732 16584
rect 32680 16541 32689 16575
rect 32689 16541 32723 16575
rect 32723 16541 32732 16575
rect 32680 16532 32732 16541
rect 33416 16600 33468 16652
rect 33232 16575 33284 16584
rect 33232 16541 33241 16575
rect 33241 16541 33275 16575
rect 33275 16541 33284 16575
rect 34060 16600 34112 16652
rect 33232 16532 33284 16541
rect 23112 16464 23164 16516
rect 24492 16464 24544 16516
rect 27068 16464 27120 16516
rect 28632 16464 28684 16516
rect 31852 16464 31904 16516
rect 36176 16532 36228 16584
rect 36912 16575 36964 16584
rect 36912 16541 36921 16575
rect 36921 16541 36955 16575
rect 36955 16541 36964 16575
rect 36912 16532 36964 16541
rect 35440 16464 35492 16516
rect 28724 16396 28776 16448
rect 30104 16396 30156 16448
rect 30472 16396 30524 16448
rect 33324 16396 33376 16448
rect 37096 16439 37148 16448
rect 37096 16405 37105 16439
rect 37105 16405 37139 16439
rect 37139 16405 37148 16439
rect 37096 16396 37148 16405
rect 4874 16294 4926 16346
rect 4938 16294 4990 16346
rect 5002 16294 5054 16346
rect 5066 16294 5118 16346
rect 5130 16294 5182 16346
rect 35594 16294 35646 16346
rect 35658 16294 35710 16346
rect 35722 16294 35774 16346
rect 35786 16294 35838 16346
rect 35850 16294 35902 16346
rect 1952 16192 2004 16244
rect 6920 16235 6972 16244
rect 6920 16201 6929 16235
rect 6929 16201 6963 16235
rect 6963 16201 6972 16235
rect 6920 16192 6972 16201
rect 9404 16192 9456 16244
rect 10140 16192 10192 16244
rect 9956 16124 10008 16176
rect 7840 16056 7892 16108
rect 7196 16031 7248 16040
rect 7196 15997 7205 16031
rect 7205 15997 7239 16031
rect 7239 15997 7248 16031
rect 7196 15988 7248 15997
rect 5540 15852 5592 15904
rect 9220 16056 9272 16108
rect 10784 16056 10836 16108
rect 12256 16192 12308 16244
rect 13820 16192 13872 16244
rect 13544 16167 13596 16176
rect 13544 16133 13553 16167
rect 13553 16133 13587 16167
rect 13587 16133 13596 16167
rect 13544 16124 13596 16133
rect 15108 16124 15160 16176
rect 15568 16192 15620 16244
rect 17132 16235 17184 16244
rect 17132 16201 17141 16235
rect 17141 16201 17175 16235
rect 17175 16201 17184 16235
rect 17132 16192 17184 16201
rect 18144 16192 18196 16244
rect 19340 16192 19392 16244
rect 20168 16192 20220 16244
rect 20444 16192 20496 16244
rect 24584 16235 24636 16244
rect 24584 16201 24593 16235
rect 24593 16201 24627 16235
rect 24627 16201 24636 16235
rect 24584 16192 24636 16201
rect 12440 16056 12492 16108
rect 12992 16056 13044 16108
rect 16948 16099 17000 16108
rect 16948 16065 16957 16099
rect 16957 16065 16991 16099
rect 16991 16065 17000 16099
rect 16948 16056 17000 16065
rect 18236 16124 18288 16176
rect 23480 16167 23532 16176
rect 18880 16099 18932 16108
rect 18880 16065 18889 16099
rect 18889 16065 18923 16099
rect 18923 16065 18932 16099
rect 18880 16056 18932 16065
rect 23480 16133 23489 16167
rect 23489 16133 23523 16167
rect 23523 16133 23532 16167
rect 23480 16124 23532 16133
rect 28632 16167 28684 16176
rect 28632 16133 28641 16167
rect 28641 16133 28675 16167
rect 28675 16133 28684 16167
rect 28632 16124 28684 16133
rect 28816 16192 28868 16244
rect 30012 16235 30064 16244
rect 30012 16201 30021 16235
rect 30021 16201 30055 16235
rect 30055 16201 30064 16235
rect 30012 16192 30064 16201
rect 9128 16031 9180 16040
rect 9128 15997 9137 16031
rect 9137 15997 9171 16031
rect 9171 15997 9180 16031
rect 9128 15988 9180 15997
rect 9588 15988 9640 16040
rect 13084 15988 13136 16040
rect 13268 16031 13320 16040
rect 13268 15997 13277 16031
rect 13277 15997 13311 16031
rect 13311 15997 13320 16031
rect 13268 15988 13320 15997
rect 14096 15988 14148 16040
rect 17960 15988 18012 16040
rect 15200 15920 15252 15972
rect 25596 16056 25648 16108
rect 27160 16056 27212 16108
rect 27712 16056 27764 16108
rect 28448 16099 28500 16108
rect 28448 16065 28458 16099
rect 28458 16065 28492 16099
rect 28492 16065 28500 16099
rect 28448 16056 28500 16065
rect 29460 16099 29512 16108
rect 29460 16065 29469 16099
rect 29469 16065 29503 16099
rect 29503 16065 29512 16099
rect 29460 16056 29512 16065
rect 29552 16099 29604 16108
rect 29552 16065 29561 16099
rect 29561 16065 29595 16099
rect 29595 16065 29604 16099
rect 29552 16056 29604 16065
rect 23388 15988 23440 16040
rect 24768 16031 24820 16040
rect 24768 15997 24777 16031
rect 24777 15997 24811 16031
rect 24811 15997 24820 16031
rect 24768 15988 24820 15997
rect 25504 16031 25556 16040
rect 25504 15997 25513 16031
rect 25513 15997 25547 16031
rect 25547 15997 25556 16031
rect 25504 15988 25556 15997
rect 28632 15988 28684 16040
rect 9036 15852 9088 15904
rect 9404 15852 9456 15904
rect 11152 15895 11204 15904
rect 11152 15861 11161 15895
rect 11161 15861 11195 15895
rect 11195 15861 11204 15895
rect 11152 15852 11204 15861
rect 21916 15852 21968 15904
rect 28540 15920 28592 15972
rect 28724 15920 28776 15972
rect 30472 16056 30524 16108
rect 32772 16124 32824 16176
rect 30932 16056 30984 16108
rect 31484 16099 31536 16108
rect 31484 16065 31493 16099
rect 31493 16065 31527 16099
rect 31527 16065 31536 16099
rect 31484 16056 31536 16065
rect 32496 16056 32548 16108
rect 32680 16099 32732 16108
rect 32680 16065 32689 16099
rect 32689 16065 32723 16099
rect 32723 16065 32732 16099
rect 35440 16124 35492 16176
rect 32680 16056 32732 16065
rect 35348 16099 35400 16108
rect 35348 16065 35357 16099
rect 35357 16065 35391 16099
rect 35391 16065 35400 16099
rect 35348 16056 35400 16065
rect 36176 16099 36228 16108
rect 34520 16031 34572 16040
rect 30748 15920 30800 15972
rect 34520 15997 34529 16031
rect 34529 15997 34563 16031
rect 34563 15997 34572 16031
rect 36176 16065 36185 16099
rect 36185 16065 36219 16099
rect 36219 16065 36228 16099
rect 36176 16056 36228 16065
rect 34520 15988 34572 15997
rect 34612 15920 34664 15972
rect 23112 15852 23164 15904
rect 26608 15852 26660 15904
rect 29000 15895 29052 15904
rect 29000 15861 29009 15895
rect 29009 15861 29043 15895
rect 29043 15861 29052 15895
rect 29000 15852 29052 15861
rect 30656 15852 30708 15904
rect 32404 15895 32456 15904
rect 32404 15861 32413 15895
rect 32413 15861 32447 15895
rect 32447 15861 32456 15895
rect 32404 15852 32456 15861
rect 34796 15852 34848 15904
rect 36084 15895 36136 15904
rect 36084 15861 36093 15895
rect 36093 15861 36127 15895
rect 36127 15861 36136 15895
rect 36084 15852 36136 15861
rect 36728 15895 36780 15904
rect 36728 15861 36737 15895
rect 36737 15861 36771 15895
rect 36771 15861 36780 15895
rect 36728 15852 36780 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 7932 15648 7984 15700
rect 11152 15648 11204 15700
rect 12992 15691 13044 15700
rect 12992 15657 13001 15691
rect 13001 15657 13035 15691
rect 13035 15657 13044 15691
rect 12992 15648 13044 15657
rect 14832 15648 14884 15700
rect 6552 15512 6604 15564
rect 8300 15512 8352 15564
rect 8944 15512 8996 15564
rect 9404 15512 9456 15564
rect 13820 15580 13872 15632
rect 23480 15648 23532 15700
rect 25504 15648 25556 15700
rect 28448 15648 28500 15700
rect 29736 15648 29788 15700
rect 23848 15580 23900 15632
rect 13268 15512 13320 15564
rect 21916 15555 21968 15564
rect 21916 15521 21925 15555
rect 21925 15521 21959 15555
rect 21959 15521 21968 15555
rect 21916 15512 21968 15521
rect 22652 15512 22704 15564
rect 5816 15487 5868 15496
rect 5816 15453 5825 15487
rect 5825 15453 5859 15487
rect 5859 15453 5868 15487
rect 5816 15444 5868 15453
rect 8484 15444 8536 15496
rect 9772 15444 9824 15496
rect 9864 15444 9916 15496
rect 6552 15419 6604 15428
rect 6552 15385 6561 15419
rect 6561 15385 6595 15419
rect 6595 15385 6604 15419
rect 6552 15376 6604 15385
rect 8392 15308 8444 15360
rect 10048 15308 10100 15360
rect 10324 15308 10376 15360
rect 15200 15444 15252 15496
rect 15384 15487 15436 15496
rect 15384 15453 15393 15487
rect 15393 15453 15427 15487
rect 15427 15453 15436 15487
rect 15384 15444 15436 15453
rect 17408 15444 17460 15496
rect 18512 15444 18564 15496
rect 21640 15487 21692 15496
rect 21640 15453 21649 15487
rect 21649 15453 21683 15487
rect 21683 15453 21692 15487
rect 21640 15444 21692 15453
rect 25872 15512 25924 15564
rect 28724 15555 28776 15564
rect 28724 15521 28733 15555
rect 28733 15521 28767 15555
rect 28767 15521 28776 15555
rect 28724 15512 28776 15521
rect 28908 15512 28960 15564
rect 32496 15648 32548 15700
rect 33324 15648 33376 15700
rect 30380 15555 30432 15564
rect 30380 15521 30389 15555
rect 30389 15521 30423 15555
rect 30423 15521 30432 15555
rect 30380 15512 30432 15521
rect 30656 15555 30708 15564
rect 30656 15521 30665 15555
rect 30665 15521 30699 15555
rect 30699 15521 30708 15555
rect 30656 15512 30708 15521
rect 34336 15555 34388 15564
rect 34336 15521 34345 15555
rect 34345 15521 34379 15555
rect 34379 15521 34388 15555
rect 34336 15512 34388 15521
rect 35624 15555 35676 15564
rect 35624 15521 35633 15555
rect 35633 15521 35667 15555
rect 35667 15521 35676 15555
rect 35624 15512 35676 15521
rect 27344 15487 27396 15496
rect 27344 15453 27353 15487
rect 27353 15453 27387 15487
rect 27387 15453 27396 15487
rect 27344 15444 27396 15453
rect 27620 15444 27672 15496
rect 28448 15487 28500 15496
rect 28448 15453 28457 15487
rect 28457 15453 28491 15487
rect 28491 15453 28500 15487
rect 28448 15444 28500 15453
rect 11980 15376 12032 15428
rect 15384 15308 15436 15360
rect 22652 15376 22704 15428
rect 26608 15376 26660 15428
rect 27068 15419 27120 15428
rect 27068 15385 27077 15419
rect 27077 15385 27111 15419
rect 27111 15385 27120 15419
rect 27068 15376 27120 15385
rect 29460 15444 29512 15496
rect 29736 15487 29788 15496
rect 29736 15453 29745 15487
rect 29745 15453 29779 15487
rect 29779 15453 29788 15487
rect 29736 15444 29788 15453
rect 30288 15444 30340 15496
rect 31760 15444 31812 15496
rect 36728 15444 36780 15496
rect 30748 15376 30800 15428
rect 33048 15376 33100 15428
rect 34060 15419 34112 15428
rect 34060 15385 34069 15419
rect 34069 15385 34103 15419
rect 34103 15385 34112 15419
rect 34060 15376 34112 15385
rect 25596 15351 25648 15360
rect 25596 15317 25605 15351
rect 25605 15317 25639 15351
rect 25639 15317 25648 15351
rect 25596 15308 25648 15317
rect 29828 15351 29880 15360
rect 29828 15317 29837 15351
rect 29837 15317 29871 15351
rect 29871 15317 29880 15351
rect 29828 15308 29880 15317
rect 30840 15308 30892 15360
rect 31484 15308 31536 15360
rect 32772 15308 32824 15360
rect 36268 15308 36320 15360
rect 4874 15206 4926 15258
rect 4938 15206 4990 15258
rect 5002 15206 5054 15258
rect 5066 15206 5118 15258
rect 5130 15206 5182 15258
rect 35594 15206 35646 15258
rect 35658 15206 35710 15258
rect 35722 15206 35774 15258
rect 35786 15206 35838 15258
rect 35850 15206 35902 15258
rect 6552 15104 6604 15156
rect 7932 15104 7984 15156
rect 8116 15104 8168 15156
rect 9128 15104 9180 15156
rect 15108 15104 15160 15156
rect 22652 15147 22704 15156
rect 22652 15113 22661 15147
rect 22661 15113 22695 15147
rect 22695 15113 22704 15147
rect 22652 15104 22704 15113
rect 27068 15104 27120 15156
rect 29552 15104 29604 15156
rect 30472 15104 30524 15156
rect 32588 15104 32640 15156
rect 33048 15104 33100 15156
rect 34336 15104 34388 15156
rect 13360 15079 13412 15088
rect 13360 15045 13369 15079
rect 13369 15045 13403 15079
rect 13403 15045 13412 15079
rect 13360 15036 13412 15045
rect 13820 15036 13872 15088
rect 14464 15079 14516 15088
rect 14464 15045 14473 15079
rect 14473 15045 14507 15079
rect 14507 15045 14516 15079
rect 14464 15036 14516 15045
rect 7012 15011 7064 15020
rect 7012 14977 7021 15011
rect 7021 14977 7055 15011
rect 7055 14977 7064 15011
rect 7012 14968 7064 14977
rect 8392 14968 8444 15020
rect 8944 15011 8996 15020
rect 8944 14977 8953 15011
rect 8953 14977 8987 15011
rect 8987 14977 8996 15011
rect 8944 14968 8996 14977
rect 10324 14968 10376 15020
rect 11704 15011 11756 15020
rect 11704 14977 11713 15011
rect 11713 14977 11747 15011
rect 11747 14977 11756 15011
rect 11704 14968 11756 14977
rect 16304 15036 16356 15088
rect 19984 15036 20036 15088
rect 26424 15036 26476 15088
rect 26516 15079 26568 15088
rect 26516 15045 26525 15079
rect 26525 15045 26559 15079
rect 26559 15045 26568 15079
rect 26516 15036 26568 15045
rect 27344 15036 27396 15088
rect 14740 15011 14792 15020
rect 14740 14977 14749 15011
rect 14749 14977 14783 15011
rect 14783 14977 14792 15011
rect 15384 15011 15436 15020
rect 14740 14968 14792 14977
rect 7196 14943 7248 14952
rect 7196 14909 7205 14943
rect 7205 14909 7239 14943
rect 7239 14909 7248 14943
rect 7196 14900 7248 14909
rect 9772 14900 9824 14952
rect 15384 14977 15393 15011
rect 15393 14977 15427 15011
rect 15427 14977 15436 15011
rect 15384 14968 15436 14977
rect 22008 14968 22060 15020
rect 24584 15011 24636 15020
rect 24584 14977 24593 15011
rect 24593 14977 24627 15011
rect 24627 14977 24636 15011
rect 24584 14968 24636 14977
rect 26700 14968 26752 15020
rect 28540 15011 28592 15020
rect 15844 14900 15896 14952
rect 22928 14900 22980 14952
rect 24032 14900 24084 14952
rect 28540 14977 28549 15011
rect 28549 14977 28583 15011
rect 28583 14977 28592 15011
rect 28540 14968 28592 14977
rect 28908 14968 28960 15020
rect 29460 15011 29512 15020
rect 29460 14977 29469 15011
rect 29469 14977 29503 15011
rect 29503 14977 29512 15011
rect 29460 14968 29512 14977
rect 30012 15036 30064 15088
rect 32128 15036 32180 15088
rect 32772 15036 32824 15088
rect 29828 15011 29880 15020
rect 29828 14977 29837 15011
rect 29837 14977 29871 15011
rect 29871 14977 29880 15011
rect 30932 15011 30984 15020
rect 29828 14968 29880 14977
rect 30932 14977 30941 15011
rect 30941 14977 30975 15011
rect 30975 14977 30984 15011
rect 30932 14968 30984 14977
rect 33324 15011 33376 15020
rect 26332 14832 26384 14884
rect 29920 14900 29972 14952
rect 28264 14832 28316 14884
rect 30840 14900 30892 14952
rect 33324 14977 33333 15011
rect 33333 14977 33367 15011
rect 33367 14977 33376 15011
rect 33324 14968 33376 14977
rect 36084 15036 36136 15088
rect 36268 15011 36320 15020
rect 36268 14977 36277 15011
rect 36277 14977 36311 15011
rect 36311 14977 36320 15011
rect 36268 14968 36320 14977
rect 32496 14900 32548 14952
rect 34244 14900 34296 14952
rect 31576 14832 31628 14884
rect 11888 14807 11940 14816
rect 11888 14773 11897 14807
rect 11897 14773 11931 14807
rect 11931 14773 11940 14807
rect 11888 14764 11940 14773
rect 12256 14764 12308 14816
rect 24768 14807 24820 14816
rect 24768 14773 24777 14807
rect 24777 14773 24811 14807
rect 24811 14773 24820 14807
rect 24768 14764 24820 14773
rect 24952 14764 25004 14816
rect 31208 14764 31260 14816
rect 32128 14764 32180 14816
rect 32496 14807 32548 14816
rect 32496 14773 32505 14807
rect 32505 14773 32539 14807
rect 32539 14773 32548 14807
rect 32496 14764 32548 14773
rect 35624 14807 35676 14816
rect 35624 14773 35633 14807
rect 35633 14773 35667 14807
rect 35667 14773 35676 14807
rect 35624 14764 35676 14773
rect 36176 14807 36228 14816
rect 36176 14773 36185 14807
rect 36185 14773 36219 14807
rect 36219 14773 36228 14807
rect 36176 14764 36228 14773
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 6920 14560 6972 14612
rect 7472 14560 7524 14612
rect 11704 14603 11756 14612
rect 11704 14569 11713 14603
rect 11713 14569 11747 14603
rect 11747 14569 11756 14603
rect 11704 14560 11756 14569
rect 24032 14560 24084 14612
rect 25596 14560 25648 14612
rect 27712 14603 27764 14612
rect 2136 14492 2188 14544
rect 6092 14467 6144 14476
rect 6092 14433 6101 14467
rect 6101 14433 6135 14467
rect 6135 14433 6144 14467
rect 6092 14424 6144 14433
rect 10968 14492 11020 14544
rect 9772 14467 9824 14476
rect 9772 14433 9781 14467
rect 9781 14433 9815 14467
rect 9815 14433 9824 14467
rect 9772 14424 9824 14433
rect 9864 14467 9916 14476
rect 9864 14433 9873 14467
rect 9873 14433 9907 14467
rect 9907 14433 9916 14467
rect 9864 14424 9916 14433
rect 10600 14424 10652 14476
rect 12256 14467 12308 14476
rect 12256 14433 12265 14467
rect 12265 14433 12299 14467
rect 12299 14433 12308 14467
rect 12256 14424 12308 14433
rect 21640 14424 21692 14476
rect 22192 14424 22244 14476
rect 22928 14467 22980 14476
rect 22928 14433 22937 14467
rect 22937 14433 22971 14467
rect 22971 14433 22980 14467
rect 22928 14424 22980 14433
rect 24860 14424 24912 14476
rect 26516 14424 26568 14476
rect 5540 14356 5592 14408
rect 8392 14399 8444 14408
rect 8392 14365 8401 14399
rect 8401 14365 8435 14399
rect 8435 14365 8444 14399
rect 8392 14356 8444 14365
rect 11244 14356 11296 14408
rect 13820 14356 13872 14408
rect 21548 14356 21600 14408
rect 23572 14399 23624 14408
rect 23572 14365 23581 14399
rect 23581 14365 23615 14399
rect 23615 14365 23624 14399
rect 23572 14356 23624 14365
rect 27712 14569 27721 14603
rect 27721 14569 27755 14603
rect 27755 14569 27764 14603
rect 27712 14560 27764 14569
rect 28448 14560 28500 14612
rect 28632 14603 28684 14612
rect 28632 14569 28641 14603
rect 28641 14569 28675 14603
rect 28675 14569 28684 14603
rect 28632 14560 28684 14569
rect 31760 14560 31812 14612
rect 34060 14560 34112 14612
rect 34244 14603 34296 14612
rect 34244 14569 34253 14603
rect 34253 14569 34287 14603
rect 34287 14569 34296 14603
rect 34244 14560 34296 14569
rect 35440 14560 35492 14612
rect 28264 14424 28316 14476
rect 28724 14492 28776 14544
rect 31208 14492 31260 14544
rect 29920 14467 29972 14476
rect 29920 14433 29929 14467
rect 29929 14433 29963 14467
rect 29963 14433 29972 14467
rect 29920 14424 29972 14433
rect 30288 14424 30340 14476
rect 7380 14288 7432 14340
rect 10692 14288 10744 14340
rect 12164 14331 12216 14340
rect 12164 14297 12173 14331
rect 12173 14297 12207 14331
rect 12207 14297 12216 14331
rect 12164 14288 12216 14297
rect 25228 14331 25280 14340
rect 8576 14263 8628 14272
rect 8576 14229 8585 14263
rect 8585 14229 8619 14263
rect 8619 14229 8628 14263
rect 8576 14220 8628 14229
rect 9312 14263 9364 14272
rect 9312 14229 9321 14263
rect 9321 14229 9355 14263
rect 9355 14229 9364 14263
rect 9312 14220 9364 14229
rect 10784 14220 10836 14272
rect 10968 14263 11020 14272
rect 10968 14229 10977 14263
rect 10977 14229 11011 14263
rect 11011 14229 11020 14263
rect 10968 14220 11020 14229
rect 13820 14220 13872 14272
rect 25228 14297 25237 14331
rect 25237 14297 25271 14331
rect 25271 14297 25280 14331
rect 25228 14288 25280 14297
rect 27252 14288 27304 14340
rect 28264 14288 28316 14340
rect 28816 14356 28868 14408
rect 29736 14356 29788 14408
rect 30012 14399 30064 14408
rect 30012 14365 30021 14399
rect 30021 14365 30055 14399
rect 30055 14365 30064 14399
rect 30012 14356 30064 14365
rect 31392 14356 31444 14408
rect 34520 14492 34572 14544
rect 35624 14492 35676 14544
rect 31576 14424 31628 14476
rect 32680 14424 32732 14476
rect 32404 14399 32456 14408
rect 32404 14365 32413 14399
rect 32413 14365 32447 14399
rect 32447 14365 32456 14399
rect 32404 14356 32456 14365
rect 33232 14356 33284 14408
rect 34796 14424 34848 14476
rect 34612 14356 34664 14408
rect 36176 14356 36228 14408
rect 33324 14288 33376 14340
rect 26700 14263 26752 14272
rect 26700 14229 26709 14263
rect 26709 14229 26743 14263
rect 26743 14229 26752 14263
rect 26700 14220 26752 14229
rect 29092 14220 29144 14272
rect 31024 14220 31076 14272
rect 33048 14263 33100 14272
rect 33048 14229 33057 14263
rect 33057 14229 33091 14263
rect 33091 14229 33100 14263
rect 33048 14220 33100 14229
rect 4874 14118 4926 14170
rect 4938 14118 4990 14170
rect 5002 14118 5054 14170
rect 5066 14118 5118 14170
rect 5130 14118 5182 14170
rect 35594 14118 35646 14170
rect 35658 14118 35710 14170
rect 35722 14118 35774 14170
rect 35786 14118 35838 14170
rect 35850 14118 35902 14170
rect 7012 14059 7064 14068
rect 7012 14025 7021 14059
rect 7021 14025 7055 14059
rect 7055 14025 7064 14059
rect 7012 14016 7064 14025
rect 7472 14059 7524 14068
rect 7472 14025 7481 14059
rect 7481 14025 7515 14059
rect 7515 14025 7524 14059
rect 7472 14016 7524 14025
rect 8300 14016 8352 14068
rect 9588 14016 9640 14068
rect 10048 14059 10100 14068
rect 10048 14025 10057 14059
rect 10057 14025 10091 14059
rect 10091 14025 10100 14059
rect 10048 14016 10100 14025
rect 10692 14016 10744 14068
rect 11060 14016 11112 14068
rect 12164 14016 12216 14068
rect 13820 14059 13872 14068
rect 13820 14025 13829 14059
rect 13829 14025 13863 14059
rect 13863 14025 13872 14059
rect 13820 14016 13872 14025
rect 21548 14016 21600 14068
rect 23480 14016 23532 14068
rect 26700 14016 26752 14068
rect 27160 14016 27212 14068
rect 30288 14059 30340 14068
rect 8576 13991 8628 14000
rect 8576 13957 8585 13991
rect 8585 13957 8619 13991
rect 8619 13957 8628 13991
rect 8576 13948 8628 13957
rect 9036 13948 9088 14000
rect 11888 13948 11940 14000
rect 13728 13948 13780 14000
rect 24032 13948 24084 14000
rect 24768 13948 24820 14000
rect 7012 13880 7064 13932
rect 8300 13923 8352 13932
rect 8300 13889 8309 13923
rect 8309 13889 8343 13923
rect 8343 13889 8352 13923
rect 8300 13880 8352 13889
rect 10508 13923 10560 13932
rect 10508 13889 10517 13923
rect 10517 13889 10551 13923
rect 10551 13889 10560 13923
rect 10508 13880 10560 13889
rect 13636 13880 13688 13932
rect 22008 13880 22060 13932
rect 24860 13923 24912 13932
rect 24860 13889 24869 13923
rect 24869 13889 24903 13923
rect 24903 13889 24912 13923
rect 24860 13880 24912 13889
rect 26976 13880 27028 13932
rect 28724 13923 28776 13932
rect 28724 13889 28733 13923
rect 28733 13889 28767 13923
rect 28767 13889 28776 13923
rect 28724 13880 28776 13889
rect 29000 13923 29052 13932
rect 9588 13812 9640 13864
rect 8208 13676 8260 13728
rect 9772 13676 9824 13728
rect 10600 13676 10652 13728
rect 13360 13812 13412 13864
rect 23572 13812 23624 13864
rect 26608 13855 26660 13864
rect 12440 13676 12492 13728
rect 23848 13744 23900 13796
rect 26608 13821 26617 13855
rect 26617 13821 26651 13855
rect 26651 13821 26660 13855
rect 26608 13812 26660 13821
rect 27436 13812 27488 13864
rect 27620 13812 27672 13864
rect 28264 13812 28316 13864
rect 29000 13889 29009 13923
rect 29009 13889 29043 13923
rect 29043 13889 29052 13923
rect 29000 13880 29052 13889
rect 29092 13923 29144 13932
rect 29092 13889 29101 13923
rect 29101 13889 29135 13923
rect 29135 13889 29144 13923
rect 29092 13880 29144 13889
rect 30288 14025 30297 14059
rect 30297 14025 30331 14059
rect 30331 14025 30340 14059
rect 30288 14016 30340 14025
rect 33232 14059 33284 14068
rect 33232 14025 33241 14059
rect 33241 14025 33275 14059
rect 33275 14025 33284 14059
rect 33232 14016 33284 14025
rect 31392 13948 31444 14000
rect 30288 13880 30340 13932
rect 30564 13880 30616 13932
rect 31484 13923 31536 13932
rect 31484 13889 31493 13923
rect 31493 13889 31527 13923
rect 31527 13889 31536 13923
rect 31484 13880 31536 13889
rect 32036 13880 32088 13932
rect 34796 13880 34848 13932
rect 32772 13855 32824 13864
rect 29184 13744 29236 13796
rect 23388 13676 23440 13728
rect 28356 13676 28408 13728
rect 31208 13744 31260 13796
rect 32128 13744 32180 13796
rect 32772 13821 32781 13855
rect 32781 13821 32815 13855
rect 32815 13821 32824 13855
rect 32772 13812 32824 13821
rect 32680 13744 32732 13796
rect 30840 13719 30892 13728
rect 30840 13685 30849 13719
rect 30849 13685 30883 13719
rect 30883 13685 30892 13719
rect 30840 13676 30892 13685
rect 31668 13719 31720 13728
rect 31668 13685 31677 13719
rect 31677 13685 31711 13719
rect 31711 13685 31720 13719
rect 31668 13676 31720 13685
rect 33784 13676 33836 13728
rect 34520 13744 34572 13796
rect 36820 13744 36872 13796
rect 37004 13676 37056 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 7380 13472 7432 13524
rect 8392 13472 8444 13524
rect 9680 13472 9732 13524
rect 12164 13472 12216 13524
rect 24584 13515 24636 13524
rect 24584 13481 24593 13515
rect 24593 13481 24627 13515
rect 24627 13481 24636 13515
rect 24584 13472 24636 13481
rect 2228 13404 2280 13456
rect 8300 13404 8352 13456
rect 9036 13404 9088 13456
rect 5816 13268 5868 13320
rect 7288 13268 7340 13320
rect 8576 13311 8628 13320
rect 8576 13277 8585 13311
rect 8585 13277 8619 13311
rect 8619 13277 8628 13311
rect 8576 13268 8628 13277
rect 9312 13268 9364 13320
rect 10048 13268 10100 13320
rect 8484 13200 8536 13252
rect 10600 13379 10652 13388
rect 10600 13345 10609 13379
rect 10609 13345 10643 13379
rect 10643 13345 10652 13379
rect 10600 13336 10652 13345
rect 12440 13268 12492 13320
rect 13820 13268 13872 13320
rect 14648 13268 14700 13320
rect 25228 13404 25280 13456
rect 23112 13379 23164 13388
rect 23112 13345 23121 13379
rect 23121 13345 23155 13379
rect 23155 13345 23164 13379
rect 23112 13336 23164 13345
rect 23388 13336 23440 13388
rect 26332 13472 26384 13524
rect 27528 13472 27580 13524
rect 28816 13472 28868 13524
rect 30472 13472 30524 13524
rect 32680 13472 32732 13524
rect 32772 13472 32824 13524
rect 33232 13472 33284 13524
rect 31208 13404 31260 13456
rect 27344 13336 27396 13388
rect 24952 13268 25004 13320
rect 10600 13200 10652 13252
rect 1584 13175 1636 13184
rect 1584 13141 1593 13175
rect 1593 13141 1627 13175
rect 1627 13141 1636 13175
rect 1584 13132 1636 13141
rect 7104 13132 7156 13184
rect 12624 13200 12676 13252
rect 26608 13268 26660 13320
rect 31944 13311 31996 13320
rect 31944 13277 31953 13311
rect 31953 13277 31987 13311
rect 31987 13277 31996 13311
rect 31944 13268 31996 13277
rect 34336 13311 34388 13320
rect 34336 13277 34345 13311
rect 34345 13277 34379 13311
rect 34379 13277 34388 13311
rect 34336 13268 34388 13277
rect 34428 13268 34480 13320
rect 13360 13132 13412 13184
rect 14188 13132 14240 13184
rect 21456 13132 21508 13184
rect 22836 13175 22888 13184
rect 22836 13141 22845 13175
rect 22845 13141 22879 13175
rect 22879 13141 22888 13175
rect 22836 13132 22888 13141
rect 22928 13175 22980 13184
rect 22928 13141 22937 13175
rect 22937 13141 22971 13175
rect 22971 13141 22980 13175
rect 22928 13132 22980 13141
rect 23664 13132 23716 13184
rect 25872 13243 25924 13252
rect 25872 13209 25881 13243
rect 25881 13209 25915 13243
rect 25915 13209 25924 13243
rect 25872 13200 25924 13209
rect 26332 13200 26384 13252
rect 26792 13200 26844 13252
rect 25044 13175 25096 13184
rect 25044 13141 25053 13175
rect 25053 13141 25087 13175
rect 25087 13141 25096 13175
rect 28816 13200 28868 13252
rect 25044 13132 25096 13141
rect 29092 13132 29144 13184
rect 31024 13200 31076 13252
rect 31668 13200 31720 13252
rect 30840 13132 30892 13184
rect 37096 13175 37148 13184
rect 37096 13141 37105 13175
rect 37105 13141 37139 13175
rect 37139 13141 37148 13175
rect 37096 13132 37148 13141
rect 4874 13030 4926 13082
rect 4938 13030 4990 13082
rect 5002 13030 5054 13082
rect 5066 13030 5118 13082
rect 5130 13030 5182 13082
rect 35594 13030 35646 13082
rect 35658 13030 35710 13082
rect 35722 13030 35774 13082
rect 35786 13030 35838 13082
rect 35850 13030 35902 13082
rect 10048 12928 10100 12980
rect 10508 12928 10560 12980
rect 10784 12971 10836 12980
rect 10784 12937 10793 12971
rect 10793 12937 10827 12971
rect 10827 12937 10836 12971
rect 10784 12928 10836 12937
rect 11060 12928 11112 12980
rect 13728 12928 13780 12980
rect 22836 12928 22888 12980
rect 23664 12971 23716 12980
rect 23664 12937 23673 12971
rect 23673 12937 23707 12971
rect 23707 12937 23716 12971
rect 23664 12928 23716 12937
rect 25872 12971 25924 12980
rect 25872 12937 25881 12971
rect 25881 12937 25915 12971
rect 25915 12937 25924 12971
rect 25872 12928 25924 12937
rect 27252 12971 27304 12980
rect 27252 12937 27261 12971
rect 27261 12937 27295 12971
rect 27295 12937 27304 12971
rect 27252 12928 27304 12937
rect 28264 12971 28316 12980
rect 28264 12937 28273 12971
rect 28273 12937 28307 12971
rect 28307 12937 28316 12971
rect 28264 12928 28316 12937
rect 28816 12971 28868 12980
rect 28816 12937 28825 12971
rect 28825 12937 28859 12971
rect 28859 12937 28868 12971
rect 28816 12928 28868 12937
rect 30564 12971 30616 12980
rect 30564 12937 30573 12971
rect 30573 12937 30607 12971
rect 30607 12937 30616 12971
rect 30564 12928 30616 12937
rect 31484 12928 31536 12980
rect 7104 12860 7156 12912
rect 8300 12860 8352 12912
rect 12808 12860 12860 12912
rect 13544 12860 13596 12912
rect 22928 12860 22980 12912
rect 25044 12860 25096 12912
rect 33232 12928 33284 12980
rect 34520 12971 34572 12980
rect 34520 12937 34529 12971
rect 34529 12937 34563 12971
rect 34563 12937 34572 12971
rect 34520 12928 34572 12937
rect 33048 12903 33100 12912
rect 33048 12869 33057 12903
rect 33057 12869 33091 12903
rect 33091 12869 33100 12903
rect 33048 12860 33100 12869
rect 33784 12860 33836 12912
rect 6092 12792 6144 12844
rect 6552 12835 6604 12844
rect 6552 12801 6561 12835
rect 6561 12801 6595 12835
rect 6595 12801 6604 12835
rect 6552 12792 6604 12801
rect 11060 12792 11112 12844
rect 12256 12792 12308 12844
rect 6828 12767 6880 12776
rect 6828 12733 6837 12767
rect 6837 12733 6871 12767
rect 6871 12733 6880 12767
rect 6828 12724 6880 12733
rect 8484 12724 8536 12776
rect 9496 12724 9548 12776
rect 9772 12767 9824 12776
rect 9772 12733 9781 12767
rect 9781 12733 9815 12767
rect 9815 12733 9824 12767
rect 9772 12724 9824 12733
rect 10600 12656 10652 12708
rect 11244 12724 11296 12776
rect 13084 12792 13136 12844
rect 13820 12792 13872 12844
rect 14464 12792 14516 12844
rect 14648 12792 14700 12844
rect 22100 12835 22152 12844
rect 22100 12801 22109 12835
rect 22109 12801 22143 12835
rect 22143 12801 22152 12835
rect 22100 12792 22152 12801
rect 22836 12792 22888 12844
rect 24032 12792 24084 12844
rect 18696 12724 18748 12776
rect 23848 12767 23900 12776
rect 23848 12733 23857 12767
rect 23857 12733 23891 12767
rect 23891 12733 23900 12767
rect 24952 12792 25004 12844
rect 23848 12724 23900 12733
rect 24584 12724 24636 12776
rect 26056 12792 26108 12844
rect 27160 12792 27212 12844
rect 27436 12792 27488 12844
rect 29000 12835 29052 12844
rect 29000 12801 29009 12835
rect 29009 12801 29043 12835
rect 29043 12801 29052 12835
rect 29000 12792 29052 12801
rect 30472 12792 30524 12844
rect 31392 12835 31444 12844
rect 31392 12801 31401 12835
rect 31401 12801 31435 12835
rect 31435 12801 31444 12835
rect 31392 12792 31444 12801
rect 31944 12792 31996 12844
rect 14188 12656 14240 12708
rect 30012 12724 30064 12776
rect 31208 12767 31260 12776
rect 31208 12733 31217 12767
rect 31217 12733 31251 12767
rect 31251 12733 31260 12767
rect 31208 12724 31260 12733
rect 31760 12656 31812 12708
rect 32128 12656 32180 12708
rect 7012 12588 7064 12640
rect 9128 12631 9180 12640
rect 9128 12597 9137 12631
rect 9137 12597 9171 12631
rect 9171 12597 9180 12631
rect 9128 12588 9180 12597
rect 11152 12588 11204 12640
rect 22376 12588 22428 12640
rect 24400 12631 24452 12640
rect 24400 12597 24409 12631
rect 24409 12597 24443 12631
rect 24443 12597 24452 12631
rect 24400 12588 24452 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 6828 12384 6880 12436
rect 8484 12384 8536 12436
rect 13544 12427 13596 12436
rect 13544 12393 13553 12427
rect 13553 12393 13587 12427
rect 13587 12393 13596 12427
rect 13544 12384 13596 12393
rect 22928 12384 22980 12436
rect 8300 12316 8352 12368
rect 9404 12316 9456 12368
rect 6552 12248 6604 12300
rect 8576 12248 8628 12300
rect 11060 12316 11112 12368
rect 24584 12316 24636 12368
rect 12440 12248 12492 12300
rect 22100 12248 22152 12300
rect 23112 12248 23164 12300
rect 24768 12248 24820 12300
rect 24860 12248 24912 12300
rect 30196 12384 30248 12436
rect 31392 12384 31444 12436
rect 28908 12316 28960 12368
rect 30656 12316 30708 12368
rect 28080 12248 28132 12300
rect 34520 12316 34572 12368
rect 32036 12291 32088 12300
rect 6184 12223 6236 12232
rect 6184 12189 6193 12223
rect 6193 12189 6227 12223
rect 6227 12189 6236 12223
rect 6184 12180 6236 12189
rect 9496 12223 9548 12232
rect 9496 12189 9505 12223
rect 9505 12189 9539 12223
rect 9539 12189 9548 12223
rect 9496 12180 9548 12189
rect 9588 12180 9640 12232
rect 11152 12223 11204 12232
rect 11152 12189 11161 12223
rect 11161 12189 11195 12223
rect 11195 12189 11204 12223
rect 11152 12180 11204 12189
rect 14464 12223 14516 12232
rect 14464 12189 14473 12223
rect 14473 12189 14507 12223
rect 14507 12189 14516 12223
rect 14464 12180 14516 12189
rect 24400 12180 24452 12232
rect 29828 12180 29880 12232
rect 29920 12223 29972 12232
rect 29920 12189 29929 12223
rect 29929 12189 29963 12223
rect 29963 12189 29972 12223
rect 32036 12257 32045 12291
rect 32045 12257 32079 12291
rect 32079 12257 32088 12291
rect 32036 12248 32088 12257
rect 29920 12180 29972 12189
rect 30932 12180 30984 12232
rect 32220 12180 32272 12232
rect 34796 12180 34848 12232
rect 7104 12155 7156 12164
rect 7104 12121 7113 12155
rect 7113 12121 7147 12155
rect 7147 12121 7156 12155
rect 7104 12112 7156 12121
rect 7840 12112 7892 12164
rect 8668 12044 8720 12096
rect 9680 12044 9732 12096
rect 10876 12044 10928 12096
rect 21456 12112 21508 12164
rect 22376 12112 22428 12164
rect 24032 12112 24084 12164
rect 27344 12112 27396 12164
rect 23296 12087 23348 12096
rect 23296 12053 23305 12087
rect 23305 12053 23339 12087
rect 23339 12053 23348 12087
rect 23296 12044 23348 12053
rect 23756 12087 23808 12096
rect 23756 12053 23765 12087
rect 23765 12053 23799 12087
rect 23799 12053 23808 12087
rect 23756 12044 23808 12053
rect 28632 12155 28684 12164
rect 28632 12121 28641 12155
rect 28641 12121 28675 12155
rect 28675 12121 28684 12155
rect 28632 12112 28684 12121
rect 33140 12155 33192 12164
rect 33140 12121 33149 12155
rect 33149 12121 33183 12155
rect 33183 12121 33192 12155
rect 33140 12112 33192 12121
rect 29552 12044 29604 12096
rect 30012 12044 30064 12096
rect 32772 12087 32824 12096
rect 32772 12053 32781 12087
rect 32781 12053 32815 12087
rect 32815 12053 32824 12087
rect 32772 12044 32824 12053
rect 33232 12087 33284 12096
rect 33232 12053 33241 12087
rect 33241 12053 33275 12087
rect 33275 12053 33284 12087
rect 33968 12087 34020 12096
rect 33232 12044 33284 12053
rect 33968 12053 33977 12087
rect 33977 12053 34011 12087
rect 34011 12053 34020 12087
rect 33968 12044 34020 12053
rect 34980 12087 35032 12096
rect 34980 12053 34989 12087
rect 34989 12053 35023 12087
rect 35023 12053 35032 12087
rect 34980 12044 35032 12053
rect 4874 11942 4926 11994
rect 4938 11942 4990 11994
rect 5002 11942 5054 11994
rect 5066 11942 5118 11994
rect 5130 11942 5182 11994
rect 35594 11942 35646 11994
rect 35658 11942 35710 11994
rect 35722 11942 35774 11994
rect 35786 11942 35838 11994
rect 35850 11942 35902 11994
rect 6184 11840 6236 11892
rect 7840 11883 7892 11892
rect 7840 11849 7849 11883
rect 7849 11849 7883 11883
rect 7883 11849 7892 11883
rect 7840 11840 7892 11849
rect 9128 11840 9180 11892
rect 9680 11840 9732 11892
rect 10232 11840 10284 11892
rect 11244 11840 11296 11892
rect 11888 11840 11940 11892
rect 24584 11883 24636 11892
rect 24584 11849 24593 11883
rect 24593 11849 24627 11883
rect 24627 11849 24636 11883
rect 24584 11840 24636 11849
rect 27344 11840 27396 11892
rect 29092 11883 29144 11892
rect 29092 11849 29101 11883
rect 29101 11849 29135 11883
rect 29135 11849 29144 11883
rect 29092 11840 29144 11849
rect 30012 11883 30064 11892
rect 30012 11849 30021 11883
rect 30021 11849 30055 11883
rect 30055 11849 30064 11883
rect 30012 11840 30064 11849
rect 32772 11840 32824 11892
rect 33232 11840 33284 11892
rect 36636 11840 36688 11892
rect 9588 11772 9640 11824
rect 13636 11772 13688 11824
rect 6920 11747 6972 11756
rect 6920 11713 6929 11747
rect 6929 11713 6963 11747
rect 6963 11713 6972 11747
rect 6920 11704 6972 11713
rect 7288 11704 7340 11756
rect 7932 11704 7984 11756
rect 7012 11679 7064 11688
rect 7012 11645 7021 11679
rect 7021 11645 7055 11679
rect 7055 11645 7064 11679
rect 7012 11636 7064 11645
rect 7196 11679 7248 11688
rect 7196 11645 7205 11679
rect 7205 11645 7239 11679
rect 7239 11645 7248 11679
rect 7196 11636 7248 11645
rect 12348 11704 12400 11756
rect 12624 11747 12676 11756
rect 12624 11713 12633 11747
rect 12633 11713 12667 11747
rect 12667 11713 12676 11747
rect 12624 11704 12676 11713
rect 14740 11704 14792 11756
rect 17868 11704 17920 11756
rect 22192 11772 22244 11824
rect 23020 11772 23072 11824
rect 24768 11772 24820 11824
rect 25320 11704 25372 11756
rect 10600 11679 10652 11688
rect 10600 11645 10609 11679
rect 10609 11645 10643 11679
rect 10643 11645 10652 11679
rect 10600 11636 10652 11645
rect 11796 11679 11848 11688
rect 11796 11645 11805 11679
rect 11805 11645 11839 11679
rect 11839 11645 11848 11679
rect 11796 11636 11848 11645
rect 22284 11679 22336 11688
rect 22284 11645 22293 11679
rect 22293 11645 22327 11679
rect 22327 11645 22336 11679
rect 22284 11636 22336 11645
rect 23756 11679 23808 11688
rect 23756 11645 23765 11679
rect 23765 11645 23799 11679
rect 23799 11645 23808 11679
rect 24676 11679 24728 11688
rect 23756 11636 23808 11645
rect 24676 11645 24685 11679
rect 24685 11645 24719 11679
rect 24719 11645 24728 11679
rect 24676 11636 24728 11645
rect 25596 11636 25648 11688
rect 26608 11772 26660 11824
rect 27528 11815 27580 11824
rect 27528 11781 27537 11815
rect 27537 11781 27571 11815
rect 27571 11781 27580 11815
rect 27528 11772 27580 11781
rect 33600 11772 33652 11824
rect 34980 11772 35032 11824
rect 26148 11704 26200 11756
rect 27620 11704 27672 11756
rect 28908 11704 28960 11756
rect 30104 11747 30156 11756
rect 30104 11713 30113 11747
rect 30113 11713 30147 11747
rect 30147 11713 30156 11747
rect 30104 11704 30156 11713
rect 30748 11704 30800 11756
rect 26240 11636 26292 11688
rect 27344 11679 27396 11688
rect 27344 11645 27353 11679
rect 27353 11645 27387 11679
rect 27387 11645 27396 11679
rect 27344 11636 27396 11645
rect 30196 11636 30248 11688
rect 31208 11679 31260 11688
rect 31208 11645 31217 11679
rect 31217 11645 31251 11679
rect 31251 11645 31260 11679
rect 31208 11636 31260 11645
rect 32036 11636 32088 11688
rect 33048 11679 33100 11688
rect 33048 11645 33057 11679
rect 33057 11645 33091 11679
rect 33091 11645 33100 11679
rect 33048 11636 33100 11645
rect 33324 11679 33376 11688
rect 33324 11645 33333 11679
rect 33333 11645 33367 11679
rect 33367 11645 33376 11679
rect 33324 11636 33376 11645
rect 29000 11568 29052 11620
rect 32220 11568 32272 11620
rect 8760 11500 8812 11552
rect 11152 11543 11204 11552
rect 11152 11509 11161 11543
rect 11161 11509 11195 11543
rect 11195 11509 11204 11543
rect 11152 11500 11204 11509
rect 23848 11500 23900 11552
rect 24308 11500 24360 11552
rect 31760 11543 31812 11552
rect 31760 11509 31769 11543
rect 31769 11509 31803 11543
rect 31803 11509 31812 11543
rect 31760 11500 31812 11509
rect 32404 11543 32456 11552
rect 32404 11509 32413 11543
rect 32413 11509 32447 11543
rect 32447 11509 32456 11543
rect 32404 11500 32456 11509
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 7104 11296 7156 11348
rect 11888 11339 11940 11348
rect 11888 11305 11897 11339
rect 11897 11305 11931 11339
rect 11931 11305 11940 11339
rect 11888 11296 11940 11305
rect 12348 11339 12400 11348
rect 12348 11305 12357 11339
rect 12357 11305 12391 11339
rect 12391 11305 12400 11339
rect 12348 11296 12400 11305
rect 22284 11339 22336 11348
rect 22284 11305 22293 11339
rect 22293 11305 22327 11339
rect 22327 11305 22336 11339
rect 22284 11296 22336 11305
rect 23020 11339 23072 11348
rect 23020 11305 23029 11339
rect 23029 11305 23063 11339
rect 23063 11305 23072 11339
rect 23020 11296 23072 11305
rect 24032 11339 24084 11348
rect 24032 11305 24041 11339
rect 24041 11305 24075 11339
rect 24075 11305 24084 11339
rect 24032 11296 24084 11305
rect 25320 11339 25372 11348
rect 25320 11305 25329 11339
rect 25329 11305 25363 11339
rect 25363 11305 25372 11339
rect 25320 11296 25372 11305
rect 30012 11296 30064 11348
rect 33968 11296 34020 11348
rect 9772 11160 9824 11212
rect 12808 11203 12860 11212
rect 12808 11169 12817 11203
rect 12817 11169 12851 11203
rect 12851 11169 12860 11203
rect 12808 11160 12860 11169
rect 6644 11092 6696 11144
rect 8668 11092 8720 11144
rect 9588 11092 9640 11144
rect 10140 11135 10192 11144
rect 10140 11101 10149 11135
rect 10149 11101 10183 11135
rect 10183 11101 10192 11135
rect 10140 11092 10192 11101
rect 14464 11092 14516 11144
rect 17224 11092 17276 11144
rect 23296 11160 23348 11212
rect 24584 11160 24636 11212
rect 24952 11228 25004 11280
rect 26608 11160 26660 11212
rect 27344 11228 27396 11280
rect 30196 11228 30248 11280
rect 33600 11228 33652 11280
rect 22836 11092 22888 11144
rect 23848 11135 23900 11144
rect 23848 11101 23857 11135
rect 23857 11101 23891 11135
rect 23891 11101 23900 11135
rect 23848 11092 23900 11101
rect 29828 11160 29880 11212
rect 33048 11160 33100 11212
rect 10416 11067 10468 11076
rect 10416 11033 10425 11067
rect 10425 11033 10459 11067
rect 10459 11033 10468 11067
rect 10416 11024 10468 11033
rect 10876 11024 10928 11076
rect 13544 11024 13596 11076
rect 24676 11024 24728 11076
rect 25596 11024 25648 11076
rect 26148 11024 26200 11076
rect 27712 11067 27764 11076
rect 6368 10999 6420 11008
rect 6368 10965 6377 10999
rect 6377 10965 6411 10999
rect 6411 10965 6420 10999
rect 6368 10956 6420 10965
rect 9496 10956 9548 11008
rect 12716 10999 12768 11008
rect 12716 10965 12725 10999
rect 12725 10965 12759 10999
rect 12759 10965 12768 10999
rect 12716 10956 12768 10965
rect 26240 10999 26292 11008
rect 26240 10965 26249 10999
rect 26249 10965 26283 10999
rect 26283 10965 26292 10999
rect 27712 11033 27721 11067
rect 27721 11033 27755 11067
rect 27755 11033 27764 11067
rect 27712 11024 27764 11033
rect 28080 11024 28132 11076
rect 34336 11092 34388 11144
rect 28908 11024 28960 11076
rect 32312 11067 32364 11076
rect 28172 10999 28224 11008
rect 26240 10956 26292 10965
rect 28172 10965 28181 10999
rect 28181 10965 28215 10999
rect 28215 10965 28224 10999
rect 28172 10956 28224 10965
rect 30932 10956 30984 11008
rect 32312 11033 32321 11067
rect 32321 11033 32355 11067
rect 32355 11033 32364 11067
rect 32312 11024 32364 11033
rect 33692 10956 33744 11008
rect 4874 10854 4926 10906
rect 4938 10854 4990 10906
rect 5002 10854 5054 10906
rect 5066 10854 5118 10906
rect 5130 10854 5182 10906
rect 35594 10854 35646 10906
rect 35658 10854 35710 10906
rect 35722 10854 35774 10906
rect 35786 10854 35838 10906
rect 35850 10854 35902 10906
rect 1860 10752 1912 10804
rect 8392 10752 8444 10804
rect 6552 10684 6604 10736
rect 10140 10752 10192 10804
rect 10232 10795 10284 10804
rect 10232 10761 10241 10795
rect 10241 10761 10275 10795
rect 10275 10761 10284 10795
rect 10232 10752 10284 10761
rect 10416 10752 10468 10804
rect 24768 10752 24820 10804
rect 26240 10752 26292 10804
rect 8760 10727 8812 10736
rect 7840 10616 7892 10668
rect 7932 10659 7984 10668
rect 7932 10625 7941 10659
rect 7941 10625 7975 10659
rect 7975 10625 7984 10659
rect 8760 10693 8769 10727
rect 8769 10693 8803 10727
rect 8803 10693 8812 10727
rect 8760 10684 8812 10693
rect 9496 10684 9548 10736
rect 11796 10684 11848 10736
rect 7932 10616 7984 10625
rect 11152 10616 11204 10668
rect 13544 10616 13596 10668
rect 17868 10659 17920 10668
rect 17868 10625 17877 10659
rect 17877 10625 17911 10659
rect 17911 10625 17920 10659
rect 17868 10616 17920 10625
rect 24308 10684 24360 10736
rect 26976 10684 27028 10736
rect 29552 10727 29604 10736
rect 29552 10693 29561 10727
rect 29561 10693 29595 10727
rect 29595 10693 29604 10727
rect 29552 10684 29604 10693
rect 30104 10752 30156 10804
rect 30472 10752 30524 10804
rect 33324 10752 33376 10804
rect 32404 10684 32456 10736
rect 33140 10684 33192 10736
rect 33600 10752 33652 10804
rect 33692 10752 33744 10804
rect 24584 10616 24636 10668
rect 26056 10616 26108 10668
rect 27068 10616 27120 10668
rect 29828 10659 29880 10668
rect 29828 10625 29837 10659
rect 29837 10625 29871 10659
rect 29871 10625 29880 10659
rect 30656 10659 30708 10668
rect 29828 10616 29880 10625
rect 30656 10625 30665 10659
rect 30665 10625 30699 10659
rect 30699 10625 30708 10659
rect 30656 10616 30708 10625
rect 31392 10616 31444 10668
rect 7012 10591 7064 10600
rect 7012 10557 7021 10591
rect 7021 10557 7055 10591
rect 7055 10557 7064 10591
rect 7012 10548 7064 10557
rect 8300 10548 8352 10600
rect 11796 10548 11848 10600
rect 18420 10548 18472 10600
rect 25964 10591 26016 10600
rect 25964 10557 25973 10591
rect 25973 10557 26007 10591
rect 26007 10557 26016 10591
rect 25964 10548 26016 10557
rect 26240 10548 26292 10600
rect 26976 10548 27028 10600
rect 28816 10548 28868 10600
rect 29460 10548 29512 10600
rect 30840 10591 30892 10600
rect 30840 10557 30849 10591
rect 30849 10557 30883 10591
rect 30883 10557 30892 10591
rect 30840 10548 30892 10557
rect 6644 10480 6696 10532
rect 33232 10616 33284 10668
rect 33692 10616 33744 10668
rect 34336 10659 34388 10668
rect 34336 10625 34345 10659
rect 34345 10625 34379 10659
rect 34379 10625 34388 10659
rect 34336 10616 34388 10625
rect 7656 10412 7708 10464
rect 13912 10455 13964 10464
rect 13912 10421 13921 10455
rect 13921 10421 13955 10455
rect 13955 10421 13964 10455
rect 13912 10412 13964 10421
rect 22560 10455 22612 10464
rect 22560 10421 22569 10455
rect 22569 10421 22603 10455
rect 22603 10421 22612 10455
rect 22560 10412 22612 10421
rect 23112 10412 23164 10464
rect 24952 10412 25004 10464
rect 30380 10412 30432 10464
rect 31852 10412 31904 10464
rect 32680 10412 32732 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 11796 10251 11848 10260
rect 11796 10217 11805 10251
rect 11805 10217 11839 10251
rect 11839 10217 11848 10251
rect 11796 10208 11848 10217
rect 25596 10208 25648 10260
rect 28632 10208 28684 10260
rect 29920 10208 29972 10260
rect 30564 10208 30616 10260
rect 31852 10208 31904 10260
rect 32312 10208 32364 10260
rect 8392 10140 8444 10192
rect 6460 10072 6512 10124
rect 25964 10140 26016 10192
rect 27712 10140 27764 10192
rect 12716 10115 12768 10124
rect 8392 10047 8444 10056
rect 8392 10013 8401 10047
rect 8401 10013 8435 10047
rect 8435 10013 8444 10047
rect 8392 10004 8444 10013
rect 12716 10081 12725 10115
rect 12725 10081 12759 10115
rect 12759 10081 12768 10115
rect 12716 10072 12768 10081
rect 15476 10072 15528 10124
rect 24584 10115 24636 10124
rect 24584 10081 24593 10115
rect 24593 10081 24627 10115
rect 24627 10081 24636 10115
rect 24584 10072 24636 10081
rect 29828 10072 29880 10124
rect 29920 10072 29972 10124
rect 30196 10072 30248 10124
rect 30840 10072 30892 10124
rect 6368 9979 6420 9988
rect 6368 9945 6377 9979
rect 6377 9945 6411 9979
rect 6411 9945 6420 9979
rect 6368 9936 6420 9945
rect 7656 9936 7708 9988
rect 7840 9911 7892 9920
rect 7840 9877 7849 9911
rect 7849 9877 7883 9911
rect 7883 9877 7892 9911
rect 7840 9868 7892 9877
rect 10784 9936 10836 9988
rect 10876 9911 10928 9920
rect 10876 9877 10885 9911
rect 10885 9877 10919 9911
rect 10919 9877 10928 9911
rect 10876 9868 10928 9877
rect 13912 10004 13964 10056
rect 23664 10004 23716 10056
rect 26424 10004 26476 10056
rect 28172 10004 28224 10056
rect 29460 10004 29512 10056
rect 31760 10004 31812 10056
rect 33600 10004 33652 10056
rect 22560 9979 22612 9988
rect 22560 9945 22569 9979
rect 22569 9945 22603 9979
rect 22603 9945 22612 9979
rect 22560 9936 22612 9945
rect 24860 9979 24912 9988
rect 24860 9945 24869 9979
rect 24869 9945 24903 9979
rect 24903 9945 24912 9979
rect 24860 9936 24912 9945
rect 25504 9936 25556 9988
rect 27436 9936 27488 9988
rect 33140 9936 33192 9988
rect 30196 9911 30248 9920
rect 30196 9877 30205 9911
rect 30205 9877 30239 9911
rect 30239 9877 30248 9911
rect 32128 9911 32180 9920
rect 30196 9868 30248 9877
rect 32128 9877 32137 9911
rect 32137 9877 32171 9911
rect 32171 9877 32180 9911
rect 32128 9868 32180 9877
rect 32956 9868 33008 9920
rect 33416 9868 33468 9920
rect 4874 9766 4926 9818
rect 4938 9766 4990 9818
rect 5002 9766 5054 9818
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 35594 9766 35646 9818
rect 35658 9766 35710 9818
rect 35722 9766 35774 9818
rect 35786 9766 35838 9818
rect 35850 9766 35902 9818
rect 8392 9664 8444 9716
rect 10232 9664 10284 9716
rect 12716 9664 12768 9716
rect 13912 9664 13964 9716
rect 10876 9596 10928 9648
rect 12072 9596 12124 9648
rect 22836 9596 22888 9648
rect 23664 9596 23716 9648
rect 27712 9664 27764 9716
rect 28816 9707 28868 9716
rect 28816 9673 28825 9707
rect 28825 9673 28859 9707
rect 28859 9673 28868 9707
rect 28816 9664 28868 9673
rect 25504 9639 25556 9648
rect 7104 9528 7156 9580
rect 7840 9528 7892 9580
rect 8300 9528 8352 9580
rect 10968 9571 11020 9580
rect 7656 9503 7708 9512
rect 7656 9469 7665 9503
rect 7665 9469 7699 9503
rect 7699 9469 7708 9503
rect 7656 9460 7708 9469
rect 8208 9460 8260 9512
rect 10968 9537 10977 9571
rect 10977 9537 11011 9571
rect 11011 9537 11020 9571
rect 10968 9528 11020 9537
rect 11704 9571 11756 9580
rect 11704 9537 11713 9571
rect 11713 9537 11747 9571
rect 11747 9537 11756 9571
rect 11704 9528 11756 9537
rect 14280 9571 14332 9580
rect 14280 9537 14289 9571
rect 14289 9537 14323 9571
rect 14323 9537 14332 9571
rect 14280 9528 14332 9537
rect 6920 9392 6972 9444
rect 9772 9392 9824 9444
rect 15108 9460 15160 9512
rect 22836 9503 22888 9512
rect 22836 9469 22845 9503
rect 22845 9469 22879 9503
rect 22879 9469 22888 9503
rect 22836 9460 22888 9469
rect 24952 9571 25004 9580
rect 24952 9537 24961 9571
rect 24961 9537 24995 9571
rect 24995 9537 25004 9571
rect 24952 9528 25004 9537
rect 25504 9605 25513 9639
rect 25513 9605 25547 9639
rect 25547 9605 25556 9639
rect 25504 9596 25556 9605
rect 27620 9639 27672 9648
rect 27620 9605 27629 9639
rect 27629 9605 27663 9639
rect 27663 9605 27672 9639
rect 27620 9596 27672 9605
rect 30196 9596 30248 9648
rect 30380 9596 30432 9648
rect 31668 9596 31720 9648
rect 33416 9596 33468 9648
rect 33876 9596 33928 9648
rect 26240 9528 26292 9580
rect 27436 9460 27488 9512
rect 24860 9392 24912 9444
rect 29828 9528 29880 9580
rect 28908 9503 28960 9512
rect 28908 9469 28917 9503
rect 28917 9469 28951 9503
rect 28951 9469 28960 9503
rect 28908 9460 28960 9469
rect 1584 9367 1636 9376
rect 1584 9333 1593 9367
rect 1593 9333 1627 9367
rect 1627 9333 1636 9367
rect 1584 9324 1636 9333
rect 9864 9324 9916 9376
rect 13912 9367 13964 9376
rect 13912 9333 13921 9367
rect 13921 9333 13955 9367
rect 13955 9333 13964 9367
rect 13912 9324 13964 9333
rect 26056 9324 26108 9376
rect 26332 9324 26384 9376
rect 34428 9528 34480 9580
rect 31760 9460 31812 9512
rect 31852 9324 31904 9376
rect 32956 9324 33008 9376
rect 36912 9460 36964 9512
rect 36912 9367 36964 9376
rect 36912 9333 36921 9367
rect 36921 9333 36955 9367
rect 36955 9333 36964 9367
rect 36912 9324 36964 9333
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 7932 9120 7984 9172
rect 10784 9163 10836 9172
rect 8116 9052 8168 9104
rect 7196 8984 7248 9036
rect 7656 8984 7708 9036
rect 7932 8916 7984 8968
rect 8208 8959 8260 8968
rect 8208 8925 8217 8959
rect 8217 8925 8251 8959
rect 8251 8925 8260 8959
rect 8208 8916 8260 8925
rect 9864 8959 9916 8968
rect 9864 8925 9873 8959
rect 9873 8925 9907 8959
rect 9907 8925 9916 8959
rect 9864 8916 9916 8925
rect 10784 9129 10793 9163
rect 10793 9129 10827 9163
rect 10827 9129 10836 9163
rect 10784 9120 10836 9129
rect 10968 9120 11020 9172
rect 27620 9120 27672 9172
rect 31392 9163 31444 9172
rect 31392 9129 31401 9163
rect 31401 9129 31435 9163
rect 31435 9129 31444 9163
rect 31392 9120 31444 9129
rect 33600 9120 33652 9172
rect 33876 9120 33928 9172
rect 14188 9052 14240 9104
rect 26240 9052 26292 9104
rect 13912 8984 13964 9036
rect 24584 8984 24636 9036
rect 25688 8984 25740 9036
rect 28356 8984 28408 9036
rect 29184 8984 29236 9036
rect 31116 8984 31168 9036
rect 32036 9027 32088 9036
rect 32036 8993 32045 9027
rect 32045 8993 32079 9027
rect 32079 8993 32088 9027
rect 32036 8984 32088 8993
rect 32496 8984 32548 9036
rect 32680 9027 32732 9036
rect 32680 8993 32689 9027
rect 32689 8993 32723 9027
rect 32723 8993 32732 9027
rect 32680 8984 32732 8993
rect 33140 8984 33192 9036
rect 13544 8959 13596 8968
rect 13544 8925 13553 8959
rect 13553 8925 13587 8959
rect 13587 8925 13596 8959
rect 13544 8916 13596 8925
rect 13636 8916 13688 8968
rect 26056 8916 26108 8968
rect 32128 8916 32180 8968
rect 32956 8959 33008 8968
rect 32956 8925 32965 8959
rect 32965 8925 32999 8959
rect 32999 8925 33008 8959
rect 32956 8916 33008 8925
rect 33784 8916 33836 8968
rect 34796 8916 34848 8968
rect 6092 8823 6144 8832
rect 6092 8789 6101 8823
rect 6101 8789 6135 8823
rect 6135 8789 6144 8823
rect 6092 8780 6144 8789
rect 7104 8780 7156 8832
rect 7380 8823 7432 8832
rect 7380 8789 7389 8823
rect 7389 8789 7423 8823
rect 7423 8789 7432 8823
rect 7380 8780 7432 8789
rect 12716 8848 12768 8900
rect 14556 8891 14608 8900
rect 14556 8857 14565 8891
rect 14565 8857 14599 8891
rect 14599 8857 14608 8891
rect 14556 8848 14608 8857
rect 24952 8891 25004 8900
rect 8024 8780 8076 8832
rect 10876 8780 10928 8832
rect 15476 8780 15528 8832
rect 16028 8823 16080 8832
rect 16028 8789 16037 8823
rect 16037 8789 16071 8823
rect 16071 8789 16080 8823
rect 16028 8780 16080 8789
rect 24952 8857 24961 8891
rect 24961 8857 24995 8891
rect 24995 8857 25004 8891
rect 24952 8848 25004 8857
rect 27160 8891 27212 8900
rect 27160 8857 27169 8891
rect 27169 8857 27203 8891
rect 27203 8857 27212 8891
rect 27160 8848 27212 8857
rect 27620 8848 27672 8900
rect 31852 8891 31904 8900
rect 31852 8857 31861 8891
rect 31861 8857 31895 8891
rect 31895 8857 31904 8891
rect 31852 8848 31904 8857
rect 33600 8848 33652 8900
rect 22284 8780 22336 8832
rect 22836 8780 22888 8832
rect 28632 8823 28684 8832
rect 28632 8789 28641 8823
rect 28641 8789 28675 8823
rect 28675 8789 28684 8823
rect 28632 8780 28684 8789
rect 4874 8678 4926 8730
rect 4938 8678 4990 8730
rect 5002 8678 5054 8730
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 35594 8678 35646 8730
rect 35658 8678 35710 8730
rect 35722 8678 35774 8730
rect 35786 8678 35838 8730
rect 35850 8678 35902 8730
rect 8208 8576 8260 8628
rect 12072 8619 12124 8628
rect 12072 8585 12081 8619
rect 12081 8585 12115 8619
rect 12115 8585 12124 8619
rect 12072 8576 12124 8585
rect 14556 8576 14608 8628
rect 15568 8576 15620 8628
rect 6092 8508 6144 8560
rect 10416 8508 10468 8560
rect 10876 8551 10928 8560
rect 10876 8517 10885 8551
rect 10885 8517 10919 8551
rect 10919 8517 10928 8551
rect 10876 8508 10928 8517
rect 5816 8483 5868 8492
rect 5816 8449 5825 8483
rect 5825 8449 5859 8483
rect 5859 8449 5868 8483
rect 5816 8440 5868 8449
rect 12440 8508 12492 8560
rect 13544 8508 13596 8560
rect 14280 8508 14332 8560
rect 14464 8483 14516 8492
rect 9220 8372 9272 8424
rect 11796 8372 11848 8424
rect 13636 8372 13688 8424
rect 7012 8304 7064 8356
rect 14464 8449 14473 8483
rect 14473 8449 14507 8483
rect 14507 8449 14516 8483
rect 14464 8440 14516 8449
rect 16028 8508 16080 8560
rect 18144 8508 18196 8560
rect 14188 8304 14240 8356
rect 14556 8304 14608 8356
rect 15476 8372 15528 8424
rect 16028 8372 16080 8424
rect 17132 8415 17184 8424
rect 17132 8381 17141 8415
rect 17141 8381 17175 8415
rect 17175 8381 17184 8415
rect 17132 8372 17184 8381
rect 26424 8576 26476 8628
rect 27620 8576 27672 8628
rect 28632 8576 28684 8628
rect 30656 8576 30708 8628
rect 31668 8619 31720 8628
rect 31668 8585 31677 8619
rect 31677 8585 31711 8619
rect 31711 8585 31720 8619
rect 31668 8576 31720 8585
rect 33600 8576 33652 8628
rect 34336 8576 34388 8628
rect 25688 8440 25740 8492
rect 26056 8440 26108 8492
rect 27804 8440 27856 8492
rect 27988 8440 28040 8492
rect 30288 8508 30340 8560
rect 30840 8508 30892 8560
rect 31116 8483 31168 8492
rect 31116 8449 31125 8483
rect 31125 8449 31159 8483
rect 31159 8449 31168 8483
rect 31116 8440 31168 8449
rect 32864 8440 32916 8492
rect 32496 8415 32548 8424
rect 21456 8304 21508 8356
rect 28724 8304 28776 8356
rect 32496 8381 32505 8415
rect 32505 8381 32539 8415
rect 32539 8381 32548 8415
rect 32496 8372 32548 8381
rect 32772 8372 32824 8424
rect 34796 8440 34848 8492
rect 34612 8304 34664 8356
rect 34796 8347 34848 8356
rect 34796 8313 34805 8347
rect 34805 8313 34839 8347
rect 34839 8313 34848 8347
rect 34796 8304 34848 8313
rect 16304 8236 16356 8288
rect 28816 8236 28868 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 5816 8032 5868 8084
rect 10416 8032 10468 8084
rect 14464 8032 14516 8084
rect 17132 8032 17184 8084
rect 18144 8032 18196 8084
rect 24952 8032 25004 8084
rect 27160 8075 27212 8084
rect 27160 8041 27169 8075
rect 27169 8041 27203 8075
rect 27203 8041 27212 8075
rect 27160 8032 27212 8041
rect 31116 8032 31168 8084
rect 15200 7964 15252 8016
rect 15384 7964 15436 8016
rect 7104 7896 7156 7948
rect 8300 7896 8352 7948
rect 13636 7939 13688 7948
rect 13636 7905 13645 7939
rect 13645 7905 13679 7939
rect 13679 7905 13688 7939
rect 13636 7896 13688 7905
rect 15568 7939 15620 7948
rect 15568 7905 15577 7939
rect 15577 7905 15611 7939
rect 15611 7905 15620 7939
rect 15568 7896 15620 7905
rect 7380 7828 7432 7880
rect 12440 7828 12492 7880
rect 13544 7828 13596 7880
rect 16304 7871 16356 7880
rect 16304 7837 16313 7871
rect 16313 7837 16347 7871
rect 16347 7837 16356 7871
rect 16304 7828 16356 7837
rect 17224 7871 17276 7880
rect 17224 7837 17233 7871
rect 17233 7837 17267 7871
rect 17267 7837 17276 7871
rect 17224 7828 17276 7837
rect 26332 7828 26384 7880
rect 30564 7964 30616 8016
rect 30932 7964 30984 8016
rect 28908 7939 28960 7948
rect 28908 7905 28917 7939
rect 28917 7905 28951 7939
rect 28951 7905 28960 7939
rect 28908 7896 28960 7905
rect 29920 7939 29972 7948
rect 29920 7905 29929 7939
rect 29929 7905 29963 7939
rect 29963 7905 29972 7939
rect 29920 7896 29972 7905
rect 28632 7828 28684 7880
rect 28816 7828 28868 7880
rect 7012 7760 7064 7812
rect 8024 7760 8076 7812
rect 12624 7760 12676 7812
rect 16212 7760 16264 7812
rect 8944 7692 8996 7744
rect 9036 7692 9088 7744
rect 14372 7735 14424 7744
rect 14372 7701 14381 7735
rect 14381 7701 14415 7735
rect 14415 7701 14424 7735
rect 14372 7692 14424 7701
rect 15476 7735 15528 7744
rect 15476 7701 15485 7735
rect 15485 7701 15519 7735
rect 15519 7701 15528 7735
rect 15476 7692 15528 7701
rect 30656 7896 30708 7948
rect 31760 7896 31812 7948
rect 33140 7896 33192 7948
rect 34336 7828 34388 7880
rect 34612 7828 34664 7880
rect 32956 7760 33008 7812
rect 32772 7735 32824 7744
rect 32772 7701 32781 7735
rect 32781 7701 32815 7735
rect 32815 7701 32824 7735
rect 32772 7692 32824 7701
rect 34152 7692 34204 7744
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 35594 7590 35646 7642
rect 35658 7590 35710 7642
rect 35722 7590 35774 7642
rect 35786 7590 35838 7642
rect 35850 7590 35902 7642
rect 7104 7488 7156 7540
rect 9036 7488 9088 7540
rect 8944 7463 8996 7472
rect 8944 7429 8953 7463
rect 8953 7429 8987 7463
rect 8987 7429 8996 7463
rect 8944 7420 8996 7429
rect 14372 7420 14424 7472
rect 9220 7395 9272 7404
rect 9220 7361 9229 7395
rect 9229 7361 9263 7395
rect 9263 7361 9272 7395
rect 9220 7352 9272 7361
rect 11796 7352 11848 7404
rect 12348 7395 12400 7404
rect 12348 7361 12357 7395
rect 12357 7361 12391 7395
rect 12391 7361 12400 7395
rect 12348 7352 12400 7361
rect 12440 7352 12492 7404
rect 15936 7395 15988 7404
rect 15936 7361 15945 7395
rect 15945 7361 15979 7395
rect 15979 7361 15988 7395
rect 15936 7352 15988 7361
rect 27344 7395 27396 7404
rect 27344 7361 27353 7395
rect 27353 7361 27387 7395
rect 27387 7361 27396 7395
rect 27344 7352 27396 7361
rect 30012 7420 30064 7472
rect 30288 7488 30340 7540
rect 30380 7420 30432 7472
rect 33692 7488 33744 7540
rect 34336 7488 34388 7540
rect 34796 7420 34848 7472
rect 15292 7327 15344 7336
rect 15292 7293 15301 7327
rect 15301 7293 15335 7327
rect 15335 7293 15344 7327
rect 15292 7284 15344 7293
rect 16028 7284 16080 7336
rect 30472 7327 30524 7336
rect 30472 7293 30481 7327
rect 30481 7293 30515 7327
rect 30515 7293 30524 7327
rect 30472 7284 30524 7293
rect 12164 7191 12216 7200
rect 12164 7157 12173 7191
rect 12173 7157 12207 7191
rect 12207 7157 12216 7191
rect 12164 7148 12216 7157
rect 12808 7148 12860 7200
rect 15476 7148 15528 7200
rect 27160 7191 27212 7200
rect 27160 7157 27169 7191
rect 27169 7157 27203 7191
rect 27203 7157 27212 7191
rect 27160 7148 27212 7157
rect 27896 7191 27948 7200
rect 27896 7157 27905 7191
rect 27905 7157 27939 7191
rect 27939 7157 27948 7191
rect 27896 7148 27948 7157
rect 29000 7191 29052 7200
rect 29000 7157 29009 7191
rect 29009 7157 29043 7191
rect 29043 7157 29052 7191
rect 29000 7148 29052 7157
rect 30288 7148 30340 7200
rect 31852 7284 31904 7336
rect 32680 7284 32732 7336
rect 33048 7327 33100 7336
rect 33048 7293 33057 7327
rect 33057 7293 33091 7327
rect 33091 7293 33100 7327
rect 33048 7284 33100 7293
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 12164 6944 12216 6996
rect 27160 6944 27212 6996
rect 28724 6944 28776 6996
rect 30840 6944 30892 6996
rect 31668 6944 31720 6996
rect 15292 6808 15344 6860
rect 28724 6808 28776 6860
rect 29828 6851 29880 6860
rect 29828 6817 29837 6851
rect 29837 6817 29871 6851
rect 29871 6817 29880 6851
rect 29828 6808 29880 6817
rect 31024 6808 31076 6860
rect 31208 6808 31260 6860
rect 31668 6808 31720 6860
rect 32956 6808 33008 6860
rect 11336 6740 11388 6792
rect 11796 6783 11848 6792
rect 11796 6749 11805 6783
rect 11805 6749 11839 6783
rect 11839 6749 11848 6783
rect 11796 6740 11848 6749
rect 16212 6783 16264 6792
rect 16212 6749 16221 6783
rect 16221 6749 16255 6783
rect 16255 6749 16264 6783
rect 16212 6740 16264 6749
rect 16856 6783 16908 6792
rect 16856 6749 16865 6783
rect 16865 6749 16899 6783
rect 16899 6749 16908 6783
rect 16856 6740 16908 6749
rect 26056 6740 26108 6792
rect 27804 6740 27856 6792
rect 28632 6740 28684 6792
rect 32772 6740 32824 6792
rect 32864 6740 32916 6792
rect 34152 6783 34204 6792
rect 34152 6749 34161 6783
rect 34161 6749 34195 6783
rect 34195 6749 34204 6783
rect 34152 6740 34204 6749
rect 12808 6672 12860 6724
rect 27896 6672 27948 6724
rect 29000 6672 29052 6724
rect 33508 6672 33560 6724
rect 14740 6604 14792 6656
rect 16120 6604 16172 6656
rect 27804 6604 27856 6656
rect 27988 6647 28040 6656
rect 27988 6613 27997 6647
rect 27997 6613 28031 6647
rect 28031 6613 28040 6647
rect 27988 6604 28040 6613
rect 28448 6647 28500 6656
rect 28448 6613 28457 6647
rect 28457 6613 28491 6647
rect 28491 6613 28500 6647
rect 28448 6604 28500 6613
rect 28908 6647 28960 6656
rect 28908 6613 28917 6647
rect 28917 6613 28951 6647
rect 28951 6613 28960 6647
rect 28908 6604 28960 6613
rect 30104 6647 30156 6656
rect 30104 6613 30113 6647
rect 30113 6613 30147 6647
rect 30147 6613 30156 6647
rect 30104 6604 30156 6613
rect 30840 6604 30892 6656
rect 31300 6647 31352 6656
rect 31300 6613 31309 6647
rect 31309 6613 31343 6647
rect 31343 6613 31352 6647
rect 31300 6604 31352 6613
rect 31576 6604 31628 6656
rect 32864 6647 32916 6656
rect 32864 6613 32873 6647
rect 32873 6613 32907 6647
rect 32907 6613 32916 6647
rect 32864 6604 32916 6613
rect 33048 6604 33100 6656
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 35594 6502 35646 6554
rect 35658 6502 35710 6554
rect 35722 6502 35774 6554
rect 35786 6502 35838 6554
rect 35850 6502 35902 6554
rect 12348 6400 12400 6452
rect 14740 6400 14792 6452
rect 16856 6400 16908 6452
rect 27344 6400 27396 6452
rect 28448 6400 28500 6452
rect 11980 6307 12032 6316
rect 11980 6273 11989 6307
rect 11989 6273 12023 6307
rect 12023 6273 12032 6307
rect 11980 6264 12032 6273
rect 12992 6307 13044 6316
rect 12992 6273 13001 6307
rect 13001 6273 13035 6307
rect 13035 6273 13044 6307
rect 12992 6264 13044 6273
rect 13268 6239 13320 6248
rect 13268 6205 13277 6239
rect 13277 6205 13311 6239
rect 13311 6205 13320 6239
rect 13268 6196 13320 6205
rect 14464 6196 14516 6248
rect 15384 6332 15436 6384
rect 17592 6332 17644 6384
rect 29092 6332 29144 6384
rect 30472 6400 30524 6452
rect 31300 6332 31352 6384
rect 33692 6332 33744 6384
rect 17316 6264 17368 6316
rect 26608 6307 26660 6316
rect 26608 6273 26617 6307
rect 26617 6273 26651 6307
rect 26651 6273 26660 6307
rect 26608 6264 26660 6273
rect 29184 6264 29236 6316
rect 30840 6264 30892 6316
rect 34244 6264 34296 6316
rect 14004 6128 14056 6180
rect 15384 6196 15436 6248
rect 15568 6239 15620 6248
rect 15568 6205 15577 6239
rect 15577 6205 15611 6239
rect 15611 6205 15620 6239
rect 15568 6196 15620 6205
rect 15752 6239 15804 6248
rect 15752 6205 15761 6239
rect 15761 6205 15795 6239
rect 15795 6205 15804 6239
rect 15752 6196 15804 6205
rect 27620 6239 27672 6248
rect 27620 6205 27629 6239
rect 27629 6205 27663 6239
rect 27663 6205 27672 6239
rect 27620 6196 27672 6205
rect 29828 6196 29880 6248
rect 30472 6239 30524 6248
rect 30472 6205 30481 6239
rect 30481 6205 30515 6239
rect 30515 6205 30524 6239
rect 30472 6196 30524 6205
rect 32680 6239 32732 6248
rect 11612 6060 11664 6112
rect 14648 6060 14700 6112
rect 16856 6060 16908 6112
rect 26332 6060 26384 6112
rect 28448 6103 28500 6112
rect 28448 6069 28457 6103
rect 28457 6069 28491 6103
rect 28491 6069 28500 6103
rect 28448 6060 28500 6069
rect 30288 6060 30340 6112
rect 32680 6205 32689 6239
rect 32689 6205 32723 6239
rect 32723 6205 32732 6239
rect 32680 6196 32732 6205
rect 33508 6060 33560 6112
rect 34428 6103 34480 6112
rect 34428 6069 34437 6103
rect 34437 6069 34471 6103
rect 34471 6069 34480 6103
rect 34428 6060 34480 6069
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 15936 5856 15988 5908
rect 27712 5856 27764 5908
rect 28908 5856 28960 5908
rect 29092 5899 29144 5908
rect 29092 5865 29101 5899
rect 29101 5865 29135 5899
rect 29135 5865 29144 5899
rect 29092 5856 29144 5865
rect 30012 5856 30064 5908
rect 34244 5856 34296 5908
rect 11612 5763 11664 5772
rect 11612 5729 11621 5763
rect 11621 5729 11655 5763
rect 11655 5729 11664 5763
rect 11612 5720 11664 5729
rect 14464 5763 14516 5772
rect 14464 5729 14473 5763
rect 14473 5729 14507 5763
rect 14507 5729 14516 5763
rect 14464 5720 14516 5729
rect 15476 5788 15528 5840
rect 15752 5788 15804 5840
rect 15292 5720 15344 5772
rect 15568 5720 15620 5772
rect 16120 5763 16172 5772
rect 16120 5729 16129 5763
rect 16129 5729 16163 5763
rect 16163 5729 16172 5763
rect 16120 5720 16172 5729
rect 26332 5763 26384 5772
rect 26332 5729 26341 5763
rect 26341 5729 26375 5763
rect 26375 5729 26384 5763
rect 26332 5720 26384 5729
rect 29736 5720 29788 5772
rect 30288 5720 30340 5772
rect 31208 5720 31260 5772
rect 7012 5652 7064 5704
rect 11336 5695 11388 5704
rect 11336 5661 11345 5695
rect 11345 5661 11379 5695
rect 11379 5661 11388 5695
rect 11336 5652 11388 5661
rect 13728 5652 13780 5704
rect 14648 5695 14700 5704
rect 14648 5661 14657 5695
rect 14657 5661 14691 5695
rect 14691 5661 14700 5695
rect 14648 5652 14700 5661
rect 25044 5652 25096 5704
rect 26056 5695 26108 5704
rect 26056 5661 26065 5695
rect 26065 5661 26099 5695
rect 26099 5661 26108 5695
rect 26056 5652 26108 5661
rect 28448 5652 28500 5704
rect 29184 5652 29236 5704
rect 30380 5652 30432 5704
rect 33508 5695 33560 5704
rect 33508 5661 33517 5695
rect 33517 5661 33551 5695
rect 33551 5661 33560 5695
rect 33508 5652 33560 5661
rect 36912 5695 36964 5704
rect 36912 5661 36921 5695
rect 36921 5661 36955 5695
rect 36955 5661 36964 5695
rect 36912 5652 36964 5661
rect 12624 5584 12676 5636
rect 1584 5559 1636 5568
rect 1584 5525 1593 5559
rect 1593 5525 1627 5559
rect 1627 5525 1636 5559
rect 1584 5516 1636 5525
rect 13084 5559 13136 5568
rect 13084 5525 13093 5559
rect 13093 5525 13127 5559
rect 13127 5525 13136 5559
rect 13084 5516 13136 5525
rect 15292 5584 15344 5636
rect 16856 5584 16908 5636
rect 31208 5627 31260 5636
rect 31208 5593 31217 5627
rect 31217 5593 31251 5627
rect 31251 5593 31260 5627
rect 31208 5584 31260 5593
rect 32588 5584 32640 5636
rect 17592 5559 17644 5568
rect 17592 5525 17601 5559
rect 17601 5525 17635 5559
rect 17635 5525 17644 5559
rect 17592 5516 17644 5525
rect 32772 5516 32824 5568
rect 37096 5559 37148 5568
rect 37096 5525 37105 5559
rect 37105 5525 37139 5559
rect 37139 5525 37148 5559
rect 37096 5516 37148 5525
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 35594 5414 35646 5466
rect 35658 5414 35710 5466
rect 35722 5414 35774 5466
rect 35786 5414 35838 5466
rect 35850 5414 35902 5466
rect 12624 5312 12676 5364
rect 12992 5312 13044 5364
rect 15292 5287 15344 5296
rect 15292 5253 15301 5287
rect 15301 5253 15335 5287
rect 15335 5253 15344 5287
rect 15292 5244 15344 5253
rect 26608 5312 26660 5364
rect 27620 5312 27672 5364
rect 30104 5312 30156 5364
rect 30472 5312 30524 5364
rect 32864 5312 32916 5364
rect 33692 5312 33744 5364
rect 12624 5176 12676 5228
rect 13084 5176 13136 5228
rect 13636 5176 13688 5228
rect 15568 5219 15620 5228
rect 15568 5185 15577 5219
rect 15577 5185 15611 5219
rect 15611 5185 15620 5219
rect 32772 5287 32824 5296
rect 32772 5253 32781 5287
rect 32781 5253 32815 5287
rect 32815 5253 32824 5287
rect 32772 5244 32824 5253
rect 15568 5176 15620 5185
rect 17040 5219 17092 5228
rect 17040 5185 17049 5219
rect 17049 5185 17083 5219
rect 17083 5185 17092 5219
rect 17040 5176 17092 5185
rect 18420 5219 18472 5228
rect 18420 5185 18429 5219
rect 18429 5185 18463 5219
rect 18463 5185 18472 5219
rect 18420 5176 18472 5185
rect 18604 5176 18656 5228
rect 27712 5176 27764 5228
rect 28540 5219 28592 5228
rect 28540 5185 28549 5219
rect 28549 5185 28583 5219
rect 28583 5185 28592 5219
rect 28540 5176 28592 5185
rect 12716 5151 12768 5160
rect 12716 5117 12725 5151
rect 12725 5117 12759 5151
rect 12759 5117 12768 5151
rect 12716 5108 12768 5117
rect 12808 5108 12860 5160
rect 29644 5151 29696 5160
rect 13544 5040 13596 5092
rect 29644 5117 29653 5151
rect 29653 5117 29687 5151
rect 29687 5117 29696 5151
rect 29644 5108 29696 5117
rect 28816 5040 28868 5092
rect 30012 5040 30064 5092
rect 10876 4972 10928 5024
rect 12072 5015 12124 5024
rect 12072 4981 12081 5015
rect 12081 4981 12115 5015
rect 12115 4981 12124 5015
rect 12072 4972 12124 4981
rect 15476 4972 15528 5024
rect 16856 5015 16908 5024
rect 16856 4981 16865 5015
rect 16865 4981 16899 5015
rect 16899 4981 16908 5015
rect 16856 4972 16908 4981
rect 18144 4972 18196 5024
rect 29000 4972 29052 5024
rect 29184 5015 29236 5024
rect 29184 4981 29193 5015
rect 29193 4981 29227 5015
rect 29227 4981 29236 5015
rect 29184 4972 29236 4981
rect 31300 5176 31352 5228
rect 31576 5176 31628 5228
rect 33784 5176 33836 5228
rect 30932 5151 30984 5160
rect 30932 5117 30941 5151
rect 30941 5117 30975 5151
rect 30975 5117 30984 5151
rect 30932 5108 30984 5117
rect 31668 5108 31720 5160
rect 32496 5108 32548 5160
rect 32864 5151 32916 5160
rect 32864 5117 32873 5151
rect 32873 5117 32907 5151
rect 32907 5117 32916 5151
rect 32864 5108 32916 5117
rect 34796 5040 34848 5092
rect 30932 4972 30984 5024
rect 32128 4972 32180 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 11980 4768 12032 4820
rect 13636 4811 13688 4820
rect 13636 4777 13645 4811
rect 13645 4777 13679 4811
rect 13679 4777 13688 4811
rect 13636 4768 13688 4777
rect 13728 4768 13780 4820
rect 18696 4768 18748 4820
rect 13268 4632 13320 4684
rect 14740 4675 14792 4684
rect 14740 4641 14749 4675
rect 14749 4641 14783 4675
rect 14783 4641 14792 4675
rect 14740 4632 14792 4641
rect 14832 4675 14884 4684
rect 14832 4641 14841 4675
rect 14841 4641 14875 4675
rect 14875 4641 14884 4675
rect 14832 4632 14884 4641
rect 15384 4632 15436 4684
rect 17408 4632 17460 4684
rect 13544 4607 13596 4616
rect 13544 4573 13553 4607
rect 13553 4573 13587 4607
rect 13587 4573 13596 4607
rect 13544 4564 13596 4573
rect 22376 4632 22428 4684
rect 19984 4607 20036 4616
rect 19984 4573 19993 4607
rect 19993 4573 20027 4607
rect 20027 4573 20036 4607
rect 19984 4564 20036 4573
rect 22652 4632 22704 4684
rect 29000 4632 29052 4684
rect 31208 4768 31260 4820
rect 32588 4768 32640 4820
rect 31484 4743 31536 4752
rect 31484 4709 31493 4743
rect 31493 4709 31527 4743
rect 31527 4709 31536 4743
rect 31484 4700 31536 4709
rect 36912 4700 36964 4752
rect 32864 4632 32916 4684
rect 12900 4496 12952 4548
rect 14556 4496 14608 4548
rect 17316 4496 17368 4548
rect 17960 4496 18012 4548
rect 10784 4428 10836 4480
rect 12348 4428 12400 4480
rect 12532 4471 12584 4480
rect 12532 4437 12541 4471
rect 12541 4437 12575 4471
rect 12575 4437 12584 4471
rect 12532 4428 12584 4437
rect 12624 4471 12676 4480
rect 12624 4437 12633 4471
rect 12633 4437 12667 4471
rect 12667 4437 12676 4471
rect 12624 4428 12676 4437
rect 12808 4428 12860 4480
rect 15936 4471 15988 4480
rect 15936 4437 15945 4471
rect 15945 4437 15979 4471
rect 15979 4437 15988 4471
rect 15936 4428 15988 4437
rect 16212 4428 16264 4480
rect 18052 4471 18104 4480
rect 18052 4437 18061 4471
rect 18061 4437 18095 4471
rect 18095 4437 18104 4471
rect 18052 4428 18104 4437
rect 18420 4471 18472 4480
rect 18420 4437 18429 4471
rect 18429 4437 18463 4471
rect 18463 4437 18472 4471
rect 18420 4428 18472 4437
rect 18604 4496 18656 4548
rect 23848 4564 23900 4616
rect 23296 4496 23348 4548
rect 18880 4428 18932 4480
rect 19616 4428 19668 4480
rect 20628 4428 20680 4480
rect 22008 4471 22060 4480
rect 22008 4437 22017 4471
rect 22017 4437 22051 4471
rect 22051 4437 22060 4471
rect 22008 4428 22060 4437
rect 22928 4471 22980 4480
rect 22928 4437 22937 4471
rect 22937 4437 22971 4471
rect 22971 4437 22980 4471
rect 22928 4428 22980 4437
rect 27528 4471 27580 4480
rect 27528 4437 27537 4471
rect 27537 4437 27571 4471
rect 27571 4437 27580 4471
rect 27528 4428 27580 4437
rect 29184 4564 29236 4616
rect 29736 4607 29788 4616
rect 29736 4573 29745 4607
rect 29745 4573 29779 4607
rect 29779 4573 29788 4607
rect 29736 4564 29788 4573
rect 32128 4607 32180 4616
rect 32128 4573 32137 4607
rect 32137 4573 32171 4607
rect 32171 4573 32180 4607
rect 32128 4564 32180 4573
rect 32772 4607 32824 4616
rect 32772 4573 32781 4607
rect 32781 4573 32815 4607
rect 32815 4573 32824 4607
rect 32772 4564 32824 4573
rect 32956 4564 33008 4616
rect 30748 4496 30800 4548
rect 28448 4428 28500 4480
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 35594 4326 35646 4378
rect 35658 4326 35710 4378
rect 35722 4326 35774 4378
rect 35786 4326 35838 4378
rect 35850 4326 35902 4378
rect 10968 4088 11020 4140
rect 12532 4224 12584 4276
rect 15660 4224 15712 4276
rect 18880 4267 18932 4276
rect 18880 4233 18889 4267
rect 18889 4233 18923 4267
rect 18923 4233 18932 4267
rect 18880 4224 18932 4233
rect 23112 4224 23164 4276
rect 14556 4156 14608 4208
rect 15476 4156 15528 4208
rect 18144 4156 18196 4208
rect 19616 4199 19668 4208
rect 19616 4165 19625 4199
rect 19625 4165 19659 4199
rect 19659 4165 19668 4199
rect 19616 4156 19668 4165
rect 20628 4156 20680 4208
rect 22008 4156 22060 4208
rect 12440 4088 12492 4140
rect 12716 4088 12768 4140
rect 16304 4131 16356 4140
rect 16304 4097 16313 4131
rect 16313 4097 16347 4131
rect 16347 4097 16356 4131
rect 16304 4088 16356 4097
rect 9864 3884 9916 3936
rect 13268 4020 13320 4072
rect 14004 4063 14056 4072
rect 12900 3952 12952 4004
rect 12624 3884 12676 3936
rect 12992 3884 13044 3936
rect 14004 4029 14013 4063
rect 14013 4029 14047 4063
rect 14047 4029 14056 4063
rect 14004 4020 14056 4029
rect 14556 4063 14608 4072
rect 14556 4029 14565 4063
rect 14565 4029 14599 4063
rect 14599 4029 14608 4063
rect 14556 4020 14608 4029
rect 16028 4063 16080 4072
rect 16028 4029 16037 4063
rect 16037 4029 16071 4063
rect 16071 4029 16080 4063
rect 16028 4020 16080 4029
rect 23388 4088 23440 4140
rect 28448 4224 28500 4276
rect 28540 4224 28592 4276
rect 29644 4224 29696 4276
rect 31484 4224 31536 4276
rect 27528 4199 27580 4208
rect 27528 4165 27537 4199
rect 27537 4165 27571 4199
rect 27571 4165 27580 4199
rect 27528 4156 27580 4165
rect 28080 4156 28132 4208
rect 17500 4020 17552 4072
rect 22008 4063 22060 4072
rect 22008 4029 22017 4063
rect 22017 4029 22051 4063
rect 22051 4029 22060 4063
rect 22008 4020 22060 4029
rect 22928 4020 22980 4072
rect 28908 4088 28960 4140
rect 23296 3952 23348 4004
rect 20628 3884 20680 3936
rect 23020 3884 23072 3936
rect 27160 3884 27212 3936
rect 28540 4020 28592 4072
rect 30012 4063 30064 4072
rect 30012 4029 30021 4063
rect 30021 4029 30055 4063
rect 30055 4029 30064 4063
rect 30748 4131 30800 4140
rect 30748 4097 30757 4131
rect 30757 4097 30791 4131
rect 30791 4097 30800 4131
rect 30748 4088 30800 4097
rect 30012 4020 30064 4029
rect 33784 4020 33836 4072
rect 29736 3952 29788 4004
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 12348 3680 12400 3732
rect 11888 3612 11940 3664
rect 12992 3612 13044 3664
rect 11336 3544 11388 3596
rect 12164 3544 12216 3596
rect 9864 3519 9916 3528
rect 9864 3485 9873 3519
rect 9873 3485 9907 3519
rect 9907 3485 9916 3519
rect 9864 3476 9916 3485
rect 12072 3476 12124 3528
rect 13084 3476 13136 3528
rect 10784 3451 10836 3460
rect 10784 3417 10793 3451
rect 10793 3417 10827 3451
rect 10827 3417 10836 3451
rect 10784 3408 10836 3417
rect 10876 3408 10928 3460
rect 12900 3408 12952 3460
rect 12348 3340 12400 3392
rect 12992 3340 13044 3392
rect 16212 3680 16264 3732
rect 17500 3723 17552 3732
rect 17500 3689 17509 3723
rect 17509 3689 17543 3723
rect 17543 3689 17552 3723
rect 17500 3680 17552 3689
rect 18420 3680 18472 3732
rect 14004 3612 14056 3664
rect 13360 3587 13412 3596
rect 13360 3553 13369 3587
rect 13369 3553 13403 3587
rect 13403 3553 13412 3587
rect 14832 3587 14884 3596
rect 13360 3544 13412 3553
rect 14832 3553 14841 3587
rect 14841 3553 14875 3587
rect 14875 3553 14884 3587
rect 14832 3544 14884 3553
rect 17040 3612 17092 3664
rect 23112 3680 23164 3732
rect 23388 3680 23440 3732
rect 28080 3723 28132 3732
rect 28080 3689 28089 3723
rect 28089 3689 28123 3723
rect 28123 3689 28132 3723
rect 28080 3680 28132 3689
rect 22008 3544 22060 3596
rect 22192 3544 22244 3596
rect 22560 3612 22612 3664
rect 23112 3587 23164 3596
rect 23112 3553 23121 3587
rect 23121 3553 23155 3587
rect 23155 3553 23164 3587
rect 23112 3544 23164 3553
rect 27160 3612 27212 3664
rect 36728 3680 36780 3732
rect 28908 3587 28960 3596
rect 14556 3476 14608 3528
rect 18052 3476 18104 3528
rect 14556 3340 14608 3392
rect 19800 3408 19852 3460
rect 19892 3408 19944 3460
rect 21916 3408 21968 3460
rect 22928 3476 22980 3528
rect 23848 3519 23900 3528
rect 23848 3485 23857 3519
rect 23857 3485 23891 3519
rect 23891 3485 23900 3519
rect 23848 3476 23900 3485
rect 24584 3476 24636 3528
rect 28908 3553 28917 3587
rect 28917 3553 28951 3587
rect 28951 3553 28960 3587
rect 28908 3544 28960 3553
rect 25044 3408 25096 3460
rect 17868 3340 17920 3392
rect 18604 3383 18656 3392
rect 18604 3349 18613 3383
rect 18613 3349 18647 3383
rect 18647 3349 18656 3383
rect 22008 3383 22060 3392
rect 18604 3340 18656 3349
rect 22008 3349 22017 3383
rect 22017 3349 22051 3383
rect 22051 3349 22060 3383
rect 22008 3340 22060 3349
rect 24676 3383 24728 3392
rect 24676 3349 24685 3383
rect 24685 3349 24719 3383
rect 24719 3349 24728 3383
rect 24676 3340 24728 3349
rect 28356 3476 28408 3528
rect 32772 3476 32824 3528
rect 28908 3340 28960 3392
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 35594 3238 35646 3290
rect 35658 3238 35710 3290
rect 35722 3238 35774 3290
rect 35786 3238 35838 3290
rect 35850 3238 35902 3290
rect 7840 3000 7892 3052
rect 12348 3068 12400 3120
rect 12992 3136 13044 3188
rect 19892 3179 19944 3188
rect 19892 3145 19901 3179
rect 19901 3145 19935 3179
rect 19935 3145 19944 3179
rect 19892 3136 19944 3145
rect 19984 3136 20036 3188
rect 21364 3136 21416 3188
rect 26240 3136 26292 3188
rect 13084 3068 13136 3120
rect 16856 3068 16908 3120
rect 18696 3068 18748 3120
rect 22192 3068 22244 3120
rect 22560 3111 22612 3120
rect 22560 3077 22569 3111
rect 22569 3077 22603 3111
rect 22603 3077 22612 3111
rect 22560 3068 22612 3077
rect 24676 3068 24728 3120
rect 1584 2839 1636 2848
rect 1584 2805 1593 2839
rect 1593 2805 1627 2839
rect 1627 2805 1636 2839
rect 1584 2796 1636 2805
rect 14924 3000 14976 3052
rect 16304 3043 16356 3052
rect 16304 3009 16313 3043
rect 16313 3009 16347 3043
rect 16347 3009 16356 3043
rect 16304 3000 16356 3009
rect 19708 3043 19760 3052
rect 19708 3009 19717 3043
rect 19717 3009 19751 3043
rect 19751 3009 19760 3043
rect 19708 3000 19760 3009
rect 19800 3000 19852 3052
rect 20536 3000 20588 3052
rect 12164 2932 12216 2984
rect 15292 2932 15344 2984
rect 17408 2975 17460 2984
rect 17408 2941 17417 2975
rect 17417 2941 17451 2975
rect 17451 2941 17460 2975
rect 17408 2932 17460 2941
rect 22652 2932 22704 2984
rect 25044 3043 25096 3052
rect 25044 3009 25053 3043
rect 25053 3009 25087 3043
rect 25087 3009 25096 3043
rect 36728 3043 36780 3052
rect 25044 3000 25096 3009
rect 36728 3009 36737 3043
rect 36737 3009 36771 3043
rect 36771 3009 36780 3043
rect 36728 3000 36780 3009
rect 24768 2975 24820 2984
rect 23020 2864 23072 2916
rect 12808 2796 12860 2848
rect 14556 2839 14608 2848
rect 14556 2805 14565 2839
rect 14565 2805 14599 2839
rect 14599 2805 14608 2839
rect 14556 2796 14608 2805
rect 18052 2796 18104 2848
rect 18604 2796 18656 2848
rect 24768 2941 24777 2975
rect 24777 2941 24811 2975
rect 24811 2941 24820 2975
rect 24768 2932 24820 2941
rect 25228 2796 25280 2848
rect 36912 2839 36964 2848
rect 36912 2805 36921 2839
rect 36921 2805 36955 2839
rect 36955 2805 36964 2839
rect 36912 2796 36964 2805
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 12440 2592 12492 2644
rect 14924 2635 14976 2644
rect 14924 2601 14933 2635
rect 14933 2601 14967 2635
rect 14967 2601 14976 2635
rect 14924 2592 14976 2601
rect 16028 2592 16080 2644
rect 17408 2592 17460 2644
rect 18696 2635 18748 2644
rect 18696 2601 18705 2635
rect 18705 2601 18739 2635
rect 18739 2601 18748 2635
rect 18696 2592 18748 2601
rect 19708 2592 19760 2644
rect 21916 2592 21968 2644
rect 24768 2635 24820 2644
rect 24768 2601 24777 2635
rect 24777 2601 24811 2635
rect 24811 2601 24820 2635
rect 24768 2592 24820 2601
rect 25228 2635 25280 2644
rect 25228 2601 25237 2635
rect 25237 2601 25271 2635
rect 25271 2601 25280 2635
rect 25228 2592 25280 2601
rect 27068 2592 27120 2644
rect 34796 2592 34848 2644
rect 10968 2524 11020 2576
rect 17592 2524 17644 2576
rect 1768 2431 1820 2440
rect 1768 2397 1777 2431
rect 1777 2397 1811 2431
rect 1811 2397 1820 2431
rect 1768 2388 1820 2397
rect 4436 2431 4488 2440
rect 4436 2397 4445 2431
rect 4445 2397 4479 2431
rect 4479 2397 4488 2431
rect 4436 2388 4488 2397
rect 7196 2431 7248 2440
rect 7196 2397 7205 2431
rect 7205 2397 7239 2431
rect 7239 2397 7248 2431
rect 7196 2388 7248 2397
rect 12164 2456 12216 2508
rect 13544 2456 13596 2508
rect 17868 2499 17920 2508
rect 11152 2431 11204 2440
rect 1400 2252 1452 2304
rect 4160 2252 4212 2304
rect 6920 2252 6972 2304
rect 9680 2295 9732 2304
rect 9680 2261 9689 2295
rect 9689 2261 9723 2295
rect 9723 2261 9732 2295
rect 9680 2252 9732 2261
rect 11152 2397 11161 2431
rect 11161 2397 11195 2431
rect 11195 2397 11204 2431
rect 11152 2388 11204 2397
rect 15936 2388 15988 2440
rect 17868 2465 17877 2499
rect 17877 2465 17911 2499
rect 17911 2465 17920 2499
rect 17868 2456 17920 2465
rect 12900 2320 12952 2372
rect 11888 2252 11940 2304
rect 17316 2388 17368 2440
rect 18052 2320 18104 2372
rect 20536 2499 20588 2508
rect 20536 2465 20545 2499
rect 20545 2465 20579 2499
rect 20579 2465 20588 2499
rect 20536 2456 20588 2465
rect 22100 2456 22152 2508
rect 21456 2431 21508 2440
rect 21456 2397 21465 2431
rect 21465 2397 21499 2431
rect 21499 2397 21508 2431
rect 21456 2388 21508 2397
rect 24584 2524 24636 2576
rect 22284 2456 22336 2508
rect 23480 2456 23532 2508
rect 23020 2388 23072 2440
rect 30196 2456 30248 2508
rect 22008 2320 22060 2372
rect 22928 2320 22980 2372
rect 17960 2252 18012 2304
rect 20444 2295 20496 2304
rect 20444 2261 20453 2295
rect 20453 2261 20487 2295
rect 20487 2261 20496 2295
rect 20444 2252 20496 2261
rect 20720 2252 20772 2304
rect 31760 2388 31812 2440
rect 34520 2388 34572 2440
rect 24492 2320 24544 2372
rect 29000 2320 29052 2372
rect 37280 2252 37332 2304
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
rect 35594 2150 35646 2202
rect 35658 2150 35710 2202
rect 35722 2150 35774 2202
rect 35786 2150 35838 2202
rect 35850 2150 35902 2202
rect 1768 2048 1820 2100
rect 20444 2048 20496 2100
rect 7196 1980 7248 2032
rect 14556 1980 14608 2032
rect 4436 1912 4488 1964
rect 18052 1912 18104 1964
rect 11152 1844 11204 1896
rect 13544 1844 13596 1896
<< metal2 >>
rect 1674 40202 1730 40893
rect 4618 40202 4674 40893
rect 7562 40202 7618 40893
rect 1674 40174 1808 40202
rect 1674 40093 1730 40174
rect 1582 38720 1638 38729
rect 1582 38655 1638 38664
rect 1596 38010 1624 38655
rect 1780 38554 1808 40174
rect 4618 40174 4752 40202
rect 4618 40093 4674 40174
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 4724 38554 4752 40174
rect 7562 40174 7696 40202
rect 7562 40093 7618 40174
rect 7668 38554 7696 40174
rect 10506 40093 10562 40893
rect 13450 40202 13506 40893
rect 16394 40202 16450 40893
rect 13096 40174 13506 40202
rect 10520 38554 10548 40093
rect 13096 38554 13124 40174
rect 13450 40093 13506 40174
rect 16316 40174 16450 40202
rect 16316 38554 16344 40174
rect 16394 40093 16450 40174
rect 19338 40093 19394 40893
rect 22282 40093 22338 40893
rect 25226 40093 25282 40893
rect 28170 40093 28226 40893
rect 31114 40093 31170 40893
rect 34058 40093 34114 40893
rect 37002 40202 37058 40893
rect 36096 40174 37058 40202
rect 1768 38548 1820 38554
rect 1768 38490 1820 38496
rect 4712 38548 4764 38554
rect 4712 38490 4764 38496
rect 7656 38548 7708 38554
rect 7656 38490 7708 38496
rect 10508 38548 10560 38554
rect 10508 38490 10560 38496
rect 13084 38548 13136 38554
rect 13084 38490 13136 38496
rect 16304 38548 16356 38554
rect 19352 38536 19380 40093
rect 22296 38554 22324 40093
rect 25240 38554 25268 40093
rect 16304 38490 16356 38496
rect 19260 38508 19380 38536
rect 22284 38548 22336 38554
rect 19064 38480 19116 38486
rect 19064 38422 19116 38428
rect 18696 38412 18748 38418
rect 18696 38354 18748 38360
rect 4804 38344 4856 38350
rect 4804 38286 4856 38292
rect 8116 38344 8168 38350
rect 8116 38286 8168 38292
rect 10140 38344 10192 38350
rect 10140 38286 10192 38292
rect 10416 38344 10468 38350
rect 10416 38286 10468 38292
rect 13084 38344 13136 38350
rect 13084 38286 13136 38292
rect 14648 38344 14700 38350
rect 14648 38286 14700 38292
rect 15016 38344 15068 38350
rect 15016 38286 15068 38292
rect 15752 38344 15804 38350
rect 15752 38286 15804 38292
rect 4816 38010 4844 38286
rect 4874 38108 5182 38117
rect 4874 38106 4880 38108
rect 4936 38106 4960 38108
rect 5016 38106 5040 38108
rect 5096 38106 5120 38108
rect 5176 38106 5182 38108
rect 4936 38054 4938 38106
rect 5118 38054 5120 38106
rect 4874 38052 4880 38054
rect 4936 38052 4960 38054
rect 5016 38052 5040 38054
rect 5096 38052 5120 38054
rect 5176 38052 5182 38054
rect 4874 38043 5182 38052
rect 8128 38010 8156 38286
rect 10152 38010 10180 38286
rect 1584 38004 1636 38010
rect 1584 37946 1636 37952
rect 4804 38004 4856 38010
rect 4804 37946 4856 37952
rect 8116 38004 8168 38010
rect 8116 37946 8168 37952
rect 10140 38004 10192 38010
rect 10140 37946 10192 37952
rect 1768 37868 1820 37874
rect 1768 37810 1820 37816
rect 8300 37868 8352 37874
rect 8300 37810 8352 37816
rect 9588 37868 9640 37874
rect 9588 37810 9640 37816
rect 10324 37868 10376 37874
rect 10324 37810 10376 37816
rect 1582 35048 1638 35057
rect 1582 34983 1638 34992
rect 1596 34950 1624 34983
rect 1584 34944 1636 34950
rect 1584 34886 1636 34892
rect 1584 31680 1636 31686
rect 1584 31622 1636 31628
rect 1596 31385 1624 31622
rect 1582 31376 1638 31385
rect 1582 31311 1638 31320
rect 1584 27872 1636 27878
rect 1584 27814 1636 27820
rect 1596 27713 1624 27814
rect 1582 27704 1638 27713
rect 1582 27639 1638 27648
rect 1584 24064 1636 24070
rect 1582 24032 1584 24041
rect 1636 24032 1638 24041
rect 1582 23967 1638 23976
rect 1582 20360 1638 20369
rect 1582 20295 1584 20304
rect 1636 20295 1638 20304
rect 1584 20266 1636 20272
rect 1780 18970 1808 37810
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 8116 37256 8168 37262
rect 8116 37198 8168 37204
rect 4874 37020 5182 37029
rect 4874 37018 4880 37020
rect 4936 37018 4960 37020
rect 5016 37018 5040 37020
rect 5096 37018 5120 37020
rect 5176 37018 5182 37020
rect 4936 36966 4938 37018
rect 5118 36966 5120 37018
rect 4874 36964 4880 36966
rect 4936 36964 4960 36966
rect 5016 36964 5040 36966
rect 5096 36964 5120 36966
rect 5176 36964 5182 36966
rect 4874 36955 5182 36964
rect 8128 36650 8156 37198
rect 8208 37188 8260 37194
rect 8208 37130 8260 37136
rect 8116 36644 8168 36650
rect 8116 36586 8168 36592
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 8024 36236 8076 36242
rect 8024 36178 8076 36184
rect 7104 36168 7156 36174
rect 7104 36110 7156 36116
rect 4874 35932 5182 35941
rect 4874 35930 4880 35932
rect 4936 35930 4960 35932
rect 5016 35930 5040 35932
rect 5096 35930 5120 35932
rect 5176 35930 5182 35932
rect 4936 35878 4938 35930
rect 5118 35878 5120 35930
rect 4874 35876 4880 35878
rect 4936 35876 4960 35878
rect 5016 35876 5040 35878
rect 5096 35876 5120 35878
rect 5176 35876 5182 35878
rect 4874 35867 5182 35876
rect 6736 35488 6788 35494
rect 6736 35430 6788 35436
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 6748 35290 6776 35430
rect 6736 35284 6788 35290
rect 6736 35226 6788 35232
rect 2044 35080 2096 35086
rect 2044 35022 2096 35028
rect 1952 31816 2004 31822
rect 1952 31758 2004 31764
rect 1860 28076 1912 28082
rect 1860 28018 1912 28024
rect 1768 18964 1820 18970
rect 1768 18906 1820 18912
rect 1584 16992 1636 16998
rect 1584 16934 1636 16940
rect 1596 16697 1624 16934
rect 1582 16688 1638 16697
rect 1582 16623 1638 16632
rect 1584 13184 1636 13190
rect 1584 13126 1636 13132
rect 1596 13025 1624 13126
rect 1582 13016 1638 13025
rect 1582 12951 1638 12960
rect 1872 10810 1900 28018
rect 1964 16250 1992 31758
rect 2056 18630 2084 35022
rect 4874 34844 5182 34853
rect 4874 34842 4880 34844
rect 4936 34842 4960 34844
rect 5016 34842 5040 34844
rect 5096 34842 5120 34844
rect 5176 34842 5182 34844
rect 4936 34790 4938 34842
rect 5118 34790 5120 34842
rect 4874 34788 4880 34790
rect 4936 34788 4960 34790
rect 5016 34788 5040 34790
rect 5096 34788 5120 34790
rect 5176 34788 5182 34790
rect 4874 34779 5182 34788
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4874 33756 5182 33765
rect 4874 33754 4880 33756
rect 4936 33754 4960 33756
rect 5016 33754 5040 33756
rect 5096 33754 5120 33756
rect 5176 33754 5182 33756
rect 4936 33702 4938 33754
rect 5118 33702 5120 33754
rect 4874 33700 4880 33702
rect 4936 33700 4960 33702
rect 5016 33700 5040 33702
rect 5096 33700 5120 33702
rect 5176 33700 5182 33702
rect 4874 33691 5182 33700
rect 6920 33584 6972 33590
rect 6920 33526 6972 33532
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 6932 33130 6960 33526
rect 7012 33312 7064 33318
rect 7012 33254 7064 33260
rect 6748 33102 6960 33130
rect 6748 32910 6776 33102
rect 7024 32978 7052 33254
rect 7012 32972 7064 32978
rect 7012 32914 7064 32920
rect 6460 32904 6512 32910
rect 6460 32846 6512 32852
rect 6736 32904 6788 32910
rect 6736 32846 6788 32852
rect 4874 32668 5182 32677
rect 4874 32666 4880 32668
rect 4936 32666 4960 32668
rect 5016 32666 5040 32668
rect 5096 32666 5120 32668
rect 5176 32666 5182 32668
rect 4936 32614 4938 32666
rect 5118 32614 5120 32666
rect 4874 32612 4880 32614
rect 4936 32612 4960 32614
rect 5016 32612 5040 32614
rect 5096 32612 5120 32614
rect 5176 32612 5182 32614
rect 4874 32603 5182 32612
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4874 31580 5182 31589
rect 4874 31578 4880 31580
rect 4936 31578 4960 31580
rect 5016 31578 5040 31580
rect 5096 31578 5120 31580
rect 5176 31578 5182 31580
rect 4936 31526 4938 31578
rect 5118 31526 5120 31578
rect 4874 31524 4880 31526
rect 4936 31524 4960 31526
rect 5016 31524 5040 31526
rect 5096 31524 5120 31526
rect 5176 31524 5182 31526
rect 4874 31515 5182 31524
rect 6472 31278 6500 32846
rect 6644 32224 6696 32230
rect 6644 32166 6696 32172
rect 6552 31680 6604 31686
rect 6552 31622 6604 31628
rect 6460 31272 6512 31278
rect 6460 31214 6512 31220
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 6472 30734 6500 31214
rect 6460 30728 6512 30734
rect 6460 30670 6512 30676
rect 4874 30492 5182 30501
rect 4874 30490 4880 30492
rect 4936 30490 4960 30492
rect 5016 30490 5040 30492
rect 5096 30490 5120 30492
rect 5176 30490 5182 30492
rect 4936 30438 4938 30490
rect 5118 30438 5120 30490
rect 4874 30436 4880 30438
rect 4936 30436 4960 30438
rect 5016 30436 5040 30438
rect 5096 30436 5120 30438
rect 5176 30436 5182 30438
rect 4874 30427 5182 30436
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 6092 29504 6144 29510
rect 6092 29446 6144 29452
rect 4874 29404 5182 29413
rect 4874 29402 4880 29404
rect 4936 29402 4960 29404
rect 5016 29402 5040 29404
rect 5096 29402 5120 29404
rect 5176 29402 5182 29404
rect 4936 29350 4938 29402
rect 5118 29350 5120 29402
rect 4874 29348 4880 29350
rect 4936 29348 4960 29350
rect 5016 29348 5040 29350
rect 5096 29348 5120 29350
rect 5176 29348 5182 29350
rect 4874 29339 5182 29348
rect 6104 29238 6132 29446
rect 6092 29232 6144 29238
rect 6092 29174 6144 29180
rect 6472 29170 6500 30670
rect 6564 30598 6592 31622
rect 6656 30666 6684 32166
rect 7116 31822 7144 36110
rect 7380 36032 7432 36038
rect 7380 35974 7432 35980
rect 7472 36032 7524 36038
rect 7472 35974 7524 35980
rect 7196 35692 7248 35698
rect 7196 35634 7248 35640
rect 7208 34746 7236 35634
rect 7392 35018 7420 35974
rect 7484 35766 7512 35974
rect 7472 35760 7524 35766
rect 7472 35702 7524 35708
rect 7380 35012 7432 35018
rect 7380 34954 7432 34960
rect 7196 34740 7248 34746
rect 7196 34682 7248 34688
rect 8036 34066 8064 36178
rect 8128 36174 8156 36586
rect 8116 36168 8168 36174
rect 8116 36110 8168 36116
rect 8116 36032 8168 36038
rect 8116 35974 8168 35980
rect 8128 35290 8156 35974
rect 8220 35766 8248 37130
rect 8312 36922 8340 37810
rect 9404 37664 9456 37670
rect 9404 37606 9456 37612
rect 9416 37330 9444 37606
rect 9404 37324 9456 37330
rect 9404 37266 9456 37272
rect 8300 36916 8352 36922
rect 8300 36858 8352 36864
rect 9404 36780 9456 36786
rect 9404 36722 9456 36728
rect 9128 36576 9180 36582
rect 9128 36518 9180 36524
rect 8300 36032 8352 36038
rect 8300 35974 8352 35980
rect 8208 35760 8260 35766
rect 8208 35702 8260 35708
rect 8116 35284 8168 35290
rect 8116 35226 8168 35232
rect 8220 35154 8248 35702
rect 8312 35494 8340 35974
rect 9140 35766 9168 36518
rect 9416 36310 9444 36722
rect 9600 36378 9628 37810
rect 10232 36848 10284 36854
rect 10232 36790 10284 36796
rect 9956 36712 10008 36718
rect 9956 36654 10008 36660
rect 9588 36372 9640 36378
rect 9588 36314 9640 36320
rect 9404 36304 9456 36310
rect 9404 36246 9456 36252
rect 9128 35760 9180 35766
rect 9128 35702 9180 35708
rect 8300 35488 8352 35494
rect 8300 35430 8352 35436
rect 8208 35148 8260 35154
rect 8208 35090 8260 35096
rect 8024 34060 8076 34066
rect 8024 34002 8076 34008
rect 7380 33856 7432 33862
rect 7380 33798 7432 33804
rect 7392 33522 7420 33798
rect 7380 33516 7432 33522
rect 7380 33458 7432 33464
rect 7288 32836 7340 32842
rect 7288 32778 7340 32784
rect 7300 32026 7328 32778
rect 7840 32360 7892 32366
rect 7840 32302 7892 32308
rect 7852 32026 7880 32302
rect 7288 32020 7340 32026
rect 7288 31962 7340 31968
rect 7840 32020 7892 32026
rect 7840 31962 7892 31968
rect 8036 31890 8064 34002
rect 8220 33998 8248 35090
rect 8852 34944 8904 34950
rect 8852 34886 8904 34892
rect 8864 34746 8892 34886
rect 8852 34740 8904 34746
rect 8852 34682 8904 34688
rect 8208 33992 8260 33998
rect 8208 33934 8260 33940
rect 8220 33590 8248 33934
rect 8484 33924 8536 33930
rect 8484 33866 8536 33872
rect 8208 33584 8260 33590
rect 8208 33526 8260 33532
rect 8392 33584 8444 33590
rect 8392 33526 8444 33532
rect 8116 33448 8168 33454
rect 8116 33390 8168 33396
rect 8128 32570 8156 33390
rect 8404 32586 8432 33526
rect 8496 33114 8524 33866
rect 9128 33856 9180 33862
rect 9128 33798 9180 33804
rect 8484 33108 8536 33114
rect 8484 33050 8536 33056
rect 8116 32564 8168 32570
rect 8116 32506 8168 32512
rect 8312 32558 8432 32586
rect 8312 32502 8340 32558
rect 8300 32496 8352 32502
rect 8300 32438 8352 32444
rect 8944 32428 8996 32434
rect 8944 32370 8996 32376
rect 8668 32224 8720 32230
rect 8668 32166 8720 32172
rect 8680 31890 8708 32166
rect 8024 31884 8076 31890
rect 8024 31826 8076 31832
rect 8668 31884 8720 31890
rect 8668 31826 8720 31832
rect 6920 31816 6972 31822
rect 6920 31758 6972 31764
rect 7104 31816 7156 31822
rect 7104 31758 7156 31764
rect 6644 30660 6696 30666
rect 6644 30602 6696 30608
rect 6552 30592 6604 30598
rect 6552 30534 6604 30540
rect 6932 29850 6960 31758
rect 7012 31340 7064 31346
rect 7012 31282 7064 31288
rect 7024 30122 7052 31282
rect 7104 30796 7156 30802
rect 7104 30738 7156 30744
rect 7012 30116 7064 30122
rect 7012 30058 7064 30064
rect 6920 29844 6972 29850
rect 6920 29786 6972 29792
rect 6932 29646 6960 29786
rect 6920 29640 6972 29646
rect 6920 29582 6972 29588
rect 6460 29164 6512 29170
rect 6460 29106 6512 29112
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 6828 28416 6880 28422
rect 6828 28358 6880 28364
rect 4874 28316 5182 28325
rect 4874 28314 4880 28316
rect 4936 28314 4960 28316
rect 5016 28314 5040 28316
rect 5096 28314 5120 28316
rect 5176 28314 5182 28316
rect 4936 28262 4938 28314
rect 5118 28262 5120 28314
rect 4874 28260 4880 28262
rect 4936 28260 4960 28262
rect 5016 28260 5040 28262
rect 5096 28260 5120 28262
rect 5176 28260 5182 28262
rect 4874 28251 5182 28260
rect 6840 28150 6868 28358
rect 7116 28218 7144 30738
rect 8036 29782 8064 31826
rect 8208 31680 8260 31686
rect 8208 31622 8260 31628
rect 8300 31680 8352 31686
rect 8300 31622 8352 31628
rect 8220 30938 8248 31622
rect 8208 30932 8260 30938
rect 8208 30874 8260 30880
rect 8220 30326 8248 30874
rect 8312 30394 8340 31622
rect 8956 31482 8984 32370
rect 9140 32366 9168 33798
rect 9416 32570 9444 36246
rect 9968 36174 9996 36654
rect 9956 36168 10008 36174
rect 9956 36110 10008 36116
rect 9968 35766 9996 36110
rect 9956 35760 10008 35766
rect 9956 35702 10008 35708
rect 9588 35488 9640 35494
rect 9588 35430 9640 35436
rect 9496 34944 9548 34950
rect 9496 34886 9548 34892
rect 9508 34066 9536 34886
rect 9600 34746 9628 35430
rect 9588 34740 9640 34746
rect 9588 34682 9640 34688
rect 9680 34468 9732 34474
rect 9680 34410 9732 34416
rect 9692 34066 9720 34410
rect 9496 34060 9548 34066
rect 9496 34002 9548 34008
rect 9680 34060 9732 34066
rect 9680 34002 9732 34008
rect 9508 33946 9536 34002
rect 9772 33992 9824 33998
rect 9508 33930 9628 33946
rect 9772 33934 9824 33940
rect 9508 33924 9640 33930
rect 9508 33918 9588 33924
rect 9588 33866 9640 33872
rect 9496 33856 9548 33862
rect 9496 33798 9548 33804
rect 9508 33114 9536 33798
rect 9600 33658 9628 33866
rect 9588 33652 9640 33658
rect 9588 33594 9640 33600
rect 9496 33108 9548 33114
rect 9496 33050 9548 33056
rect 9680 32904 9732 32910
rect 9680 32846 9732 32852
rect 9404 32564 9456 32570
rect 9404 32506 9456 32512
rect 9312 32428 9364 32434
rect 9312 32370 9364 32376
rect 9128 32360 9180 32366
rect 9128 32302 9180 32308
rect 9220 32224 9272 32230
rect 9220 32166 9272 32172
rect 9128 31816 9180 31822
rect 9128 31758 9180 31764
rect 8944 31476 8996 31482
rect 8944 31418 8996 31424
rect 8300 30388 8352 30394
rect 8300 30330 8352 30336
rect 8208 30320 8260 30326
rect 8208 30262 8260 30268
rect 8300 30252 8352 30258
rect 8300 30194 8352 30200
rect 8208 30184 8260 30190
rect 8208 30126 8260 30132
rect 8024 29776 8076 29782
rect 8024 29718 8076 29724
rect 7288 29504 7340 29510
rect 7288 29446 7340 29452
rect 8116 29504 8168 29510
rect 8116 29446 8168 29452
rect 7300 29238 7328 29446
rect 8128 29238 8156 29446
rect 7288 29232 7340 29238
rect 7288 29174 7340 29180
rect 8116 29232 8168 29238
rect 8116 29174 8168 29180
rect 8220 28626 8248 30126
rect 8312 29714 8340 30194
rect 9140 30122 9168 31758
rect 9232 31414 9260 32166
rect 9220 31408 9272 31414
rect 9220 31350 9272 31356
rect 9220 30728 9272 30734
rect 9324 30716 9352 32370
rect 9692 31770 9720 32846
rect 9784 31822 9812 33934
rect 10140 33584 10192 33590
rect 10140 33526 10192 33532
rect 10048 33516 10100 33522
rect 10048 33458 10100 33464
rect 10060 32978 10088 33458
rect 10048 32972 10100 32978
rect 10048 32914 10100 32920
rect 9600 31742 9720 31770
rect 9772 31816 9824 31822
rect 9772 31758 9824 31764
rect 9404 31136 9456 31142
rect 9404 31078 9456 31084
rect 9272 30688 9352 30716
rect 9220 30670 9272 30676
rect 9128 30116 9180 30122
rect 9128 30058 9180 30064
rect 9232 29850 9260 30670
rect 9312 30592 9364 30598
rect 9312 30534 9364 30540
rect 8760 29844 8812 29850
rect 8760 29786 8812 29792
rect 9220 29844 9272 29850
rect 9220 29786 9272 29792
rect 8300 29708 8352 29714
rect 8300 29650 8352 29656
rect 8208 28620 8260 28626
rect 8208 28562 8260 28568
rect 7104 28212 7156 28218
rect 7104 28154 7156 28160
rect 6828 28144 6880 28150
rect 6828 28086 6880 28092
rect 7288 28144 7340 28150
rect 7288 28086 7340 28092
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 7300 27606 7328 28086
rect 7288 27600 7340 27606
rect 7288 27542 7340 27548
rect 8220 27538 8248 28562
rect 8312 28422 8340 29650
rect 8392 29504 8444 29510
rect 8392 29446 8444 29452
rect 8404 28966 8432 29446
rect 8392 28960 8444 28966
rect 8392 28902 8444 28908
rect 8300 28416 8352 28422
rect 8300 28358 8352 28364
rect 8312 28218 8340 28358
rect 8300 28212 8352 28218
rect 8300 28154 8352 28160
rect 8772 28082 8800 29786
rect 9324 29306 9352 30534
rect 9416 30394 9444 31078
rect 9404 30388 9456 30394
rect 9404 30330 9456 30336
rect 9600 30190 9628 31742
rect 9784 30802 9812 31758
rect 9772 30796 9824 30802
rect 9772 30738 9824 30744
rect 9588 30184 9640 30190
rect 10152 30138 10180 33526
rect 9588 30126 9640 30132
rect 9312 29300 9364 29306
rect 9312 29242 9364 29248
rect 9312 29096 9364 29102
rect 9600 29050 9628 30126
rect 9312 29038 9364 29044
rect 9220 28416 9272 28422
rect 9220 28358 9272 28364
rect 8760 28076 8812 28082
rect 8760 28018 8812 28024
rect 8208 27532 8260 27538
rect 8208 27474 8260 27480
rect 8772 27470 8800 28018
rect 8760 27464 8812 27470
rect 8760 27406 8812 27412
rect 7932 27328 7984 27334
rect 7932 27270 7984 27276
rect 4874 27228 5182 27237
rect 4874 27226 4880 27228
rect 4936 27226 4960 27228
rect 5016 27226 5040 27228
rect 5096 27226 5120 27228
rect 5176 27226 5182 27228
rect 4936 27174 4938 27226
rect 5118 27174 5120 27226
rect 4874 27172 4880 27174
rect 4936 27172 4960 27174
rect 5016 27172 5040 27174
rect 5096 27172 5120 27174
rect 5176 27172 5182 27174
rect 4874 27163 5182 27172
rect 7748 26920 7800 26926
rect 7748 26862 7800 26868
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 7760 26586 7788 26862
rect 7748 26580 7800 26586
rect 7748 26522 7800 26528
rect 7944 26382 7972 27270
rect 8392 27056 8444 27062
rect 8392 26998 8444 27004
rect 8404 26586 8432 26998
rect 8392 26580 8444 26586
rect 8392 26522 8444 26528
rect 8772 26382 8800 27406
rect 9232 27334 9260 28358
rect 9324 28014 9352 29038
rect 9508 29022 9628 29050
rect 10060 30110 10180 30138
rect 9508 28694 9536 29022
rect 9588 28960 9640 28966
rect 9588 28902 9640 28908
rect 9496 28688 9548 28694
rect 9496 28630 9548 28636
rect 9600 28626 9628 28902
rect 9588 28620 9640 28626
rect 9588 28562 9640 28568
rect 9312 28008 9364 28014
rect 9312 27950 9364 27956
rect 9324 27538 9352 27950
rect 9312 27532 9364 27538
rect 9312 27474 9364 27480
rect 9588 27464 9640 27470
rect 9588 27406 9640 27412
rect 9220 27328 9272 27334
rect 9220 27270 9272 27276
rect 9232 27130 9260 27270
rect 9600 27130 9628 27406
rect 9680 27396 9732 27402
rect 9680 27338 9732 27344
rect 9692 27130 9720 27338
rect 9220 27124 9272 27130
rect 9220 27066 9272 27072
rect 9588 27124 9640 27130
rect 9588 27066 9640 27072
rect 9680 27124 9732 27130
rect 9680 27066 9732 27072
rect 9036 26784 9088 26790
rect 9036 26726 9088 26732
rect 7932 26376 7984 26382
rect 7932 26318 7984 26324
rect 8760 26376 8812 26382
rect 8760 26318 8812 26324
rect 9048 26234 9076 26726
rect 10060 26518 10088 30110
rect 10140 30048 10192 30054
rect 10140 29990 10192 29996
rect 10152 29646 10180 29990
rect 10140 29640 10192 29646
rect 10140 29582 10192 29588
rect 10048 26512 10100 26518
rect 10048 26454 10100 26460
rect 10060 26382 10088 26454
rect 10048 26376 10100 26382
rect 10048 26318 10100 26324
rect 9680 26240 9732 26246
rect 9048 26206 9168 26234
rect 4874 26140 5182 26149
rect 4874 26138 4880 26140
rect 4936 26138 4960 26140
rect 5016 26138 5040 26140
rect 5096 26138 5120 26140
rect 5176 26138 5182 26140
rect 4936 26086 4938 26138
rect 5118 26086 5120 26138
rect 4874 26084 4880 26086
rect 4936 26084 4960 26086
rect 5016 26084 5040 26086
rect 5096 26084 5120 26086
rect 5176 26084 5182 26086
rect 4874 26075 5182 26084
rect 9140 25906 9168 26206
rect 9680 26182 9732 26188
rect 10140 26240 10192 26246
rect 10140 26182 10192 26188
rect 9128 25900 9180 25906
rect 9128 25842 9180 25848
rect 8576 25832 8628 25838
rect 8576 25774 8628 25780
rect 8484 25696 8536 25702
rect 8484 25638 8536 25644
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 7932 25288 7984 25294
rect 7932 25230 7984 25236
rect 7748 25152 7800 25158
rect 7748 25094 7800 25100
rect 4874 25052 5182 25061
rect 4874 25050 4880 25052
rect 4936 25050 4960 25052
rect 5016 25050 5040 25052
rect 5096 25050 5120 25052
rect 5176 25050 5182 25052
rect 4936 24998 4938 25050
rect 5118 24998 5120 25050
rect 4874 24996 4880 24998
rect 4936 24996 4960 24998
rect 5016 24996 5040 24998
rect 5096 24996 5120 24998
rect 5176 24996 5182 24998
rect 4874 24987 5182 24996
rect 7760 24886 7788 25094
rect 7748 24880 7800 24886
rect 7748 24822 7800 24828
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 7944 24410 7972 25230
rect 8208 25220 8260 25226
rect 8208 25162 8260 25168
rect 7932 24404 7984 24410
rect 7932 24346 7984 24352
rect 8116 24336 8168 24342
rect 8116 24278 8168 24284
rect 2228 24200 2280 24206
rect 2228 24142 2280 24148
rect 2136 20460 2188 20466
rect 2136 20402 2188 20408
rect 2044 18624 2096 18630
rect 2044 18566 2096 18572
rect 1952 16244 2004 16250
rect 1952 16186 2004 16192
rect 2148 14550 2176 20402
rect 2136 14544 2188 14550
rect 2136 14486 2188 14492
rect 2240 13462 2268 24142
rect 7288 24064 7340 24070
rect 7288 24006 7340 24012
rect 4874 23964 5182 23973
rect 4874 23962 4880 23964
rect 4936 23962 4960 23964
rect 5016 23962 5040 23964
rect 5096 23962 5120 23964
rect 5176 23962 5182 23964
rect 4936 23910 4938 23962
rect 5118 23910 5120 23962
rect 4874 23908 4880 23910
rect 4936 23908 4960 23910
rect 5016 23908 5040 23910
rect 5096 23908 5120 23910
rect 5176 23908 5182 23910
rect 4874 23899 5182 23908
rect 7300 23798 7328 24006
rect 7288 23792 7340 23798
rect 7288 23734 7340 23740
rect 6920 23656 6972 23662
rect 6920 23598 6972 23604
rect 7288 23656 7340 23662
rect 7288 23598 7340 23604
rect 6932 23474 6960 23598
rect 6840 23446 6960 23474
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4874 22876 5182 22885
rect 4874 22874 4880 22876
rect 4936 22874 4960 22876
rect 5016 22874 5040 22876
rect 5096 22874 5120 22876
rect 5176 22874 5182 22876
rect 4936 22822 4938 22874
rect 5118 22822 5120 22874
rect 4874 22820 4880 22822
rect 4936 22820 4960 22822
rect 5016 22820 5040 22822
rect 5096 22820 5120 22822
rect 5176 22820 5182 22822
rect 4874 22811 5182 22820
rect 6840 22710 6868 23446
rect 7300 23322 7328 23598
rect 7288 23316 7340 23322
rect 7288 23258 7340 23264
rect 7564 23316 7616 23322
rect 7564 23258 7616 23264
rect 7576 23050 7604 23258
rect 8128 23186 8156 24278
rect 8220 24274 8248 25162
rect 8496 24886 8524 25638
rect 8588 25498 8616 25774
rect 8576 25492 8628 25498
rect 8576 25434 8628 25440
rect 9588 25356 9640 25362
rect 9588 25298 9640 25304
rect 9312 25152 9364 25158
rect 9312 25094 9364 25100
rect 8484 24880 8536 24886
rect 8484 24822 8536 24828
rect 9128 24608 9180 24614
rect 9128 24550 9180 24556
rect 9220 24608 9272 24614
rect 9220 24550 9272 24556
rect 9140 24274 9168 24550
rect 8208 24268 8260 24274
rect 8208 24210 8260 24216
rect 9128 24268 9180 24274
rect 9128 24210 9180 24216
rect 8116 23180 8168 23186
rect 8116 23122 8168 23128
rect 7564 23044 7616 23050
rect 7564 22986 7616 22992
rect 6920 22976 6972 22982
rect 6920 22918 6972 22924
rect 7472 22976 7524 22982
rect 7472 22918 7524 22924
rect 6932 22778 6960 22918
rect 6920 22772 6972 22778
rect 6920 22714 6972 22720
rect 6828 22704 6880 22710
rect 6828 22646 6880 22652
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4874 21788 5182 21797
rect 4874 21786 4880 21788
rect 4936 21786 4960 21788
rect 5016 21786 5040 21788
rect 5096 21786 5120 21788
rect 5176 21786 5182 21788
rect 4936 21734 4938 21786
rect 5118 21734 5120 21786
rect 4874 21732 4880 21734
rect 4936 21732 4960 21734
rect 5016 21732 5040 21734
rect 5096 21732 5120 21734
rect 5176 21732 5182 21734
rect 4874 21723 5182 21732
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 6840 21010 6868 22646
rect 6920 22568 6972 22574
rect 6920 22510 6972 22516
rect 6932 22234 6960 22510
rect 6920 22228 6972 22234
rect 6920 22170 6972 22176
rect 7484 22030 7512 22918
rect 8220 22778 8248 24210
rect 8760 23656 8812 23662
rect 8760 23598 8812 23604
rect 8576 23112 8628 23118
rect 8576 23054 8628 23060
rect 8208 22772 8260 22778
rect 8208 22714 8260 22720
rect 8024 22636 8076 22642
rect 8024 22578 8076 22584
rect 8036 22098 8064 22578
rect 8024 22092 8076 22098
rect 8024 22034 8076 22040
rect 8300 22092 8352 22098
rect 8300 22034 8352 22040
rect 7472 22024 7524 22030
rect 7472 21966 7524 21972
rect 8312 21554 8340 22034
rect 8300 21548 8352 21554
rect 8300 21490 8352 21496
rect 7840 21344 7892 21350
rect 7840 21286 7892 21292
rect 6828 21004 6880 21010
rect 6828 20946 6880 20952
rect 4874 20700 5182 20709
rect 4874 20698 4880 20700
rect 4936 20698 4960 20700
rect 5016 20698 5040 20700
rect 5096 20698 5120 20700
rect 5176 20698 5182 20700
rect 4936 20646 4938 20698
rect 5118 20646 5120 20698
rect 4874 20644 4880 20646
rect 4936 20644 4960 20646
rect 5016 20644 5040 20646
rect 5096 20644 5120 20646
rect 5176 20644 5182 20646
rect 4874 20635 5182 20644
rect 6840 20534 6868 20946
rect 7852 20874 7880 21286
rect 8588 21146 8616 23054
rect 8772 22982 8800 23598
rect 8760 22976 8812 22982
rect 8760 22918 8812 22924
rect 8576 21140 8628 21146
rect 8576 21082 8628 21088
rect 8588 21026 8616 21082
rect 8496 20998 8616 21026
rect 7104 20868 7156 20874
rect 7104 20810 7156 20816
rect 7840 20868 7892 20874
rect 7840 20810 7892 20816
rect 7116 20602 7144 20810
rect 7104 20596 7156 20602
rect 7104 20538 7156 20544
rect 6828 20528 6880 20534
rect 6828 20470 6880 20476
rect 8300 20528 8352 20534
rect 8300 20470 8352 20476
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4874 19612 5182 19621
rect 4874 19610 4880 19612
rect 4936 19610 4960 19612
rect 5016 19610 5040 19612
rect 5096 19610 5120 19612
rect 5176 19610 5182 19612
rect 4936 19558 4938 19610
rect 5118 19558 5120 19610
rect 4874 19556 4880 19558
rect 4936 19556 4960 19558
rect 5016 19556 5040 19558
rect 5096 19556 5120 19558
rect 5176 19556 5182 19558
rect 4874 19547 5182 19556
rect 8312 19446 8340 20470
rect 8496 20466 8524 20998
rect 8772 20874 8800 22918
rect 9140 22642 9168 24210
rect 9232 24138 9260 24550
rect 9220 24132 9272 24138
rect 9220 24074 9272 24080
rect 9232 22982 9260 24074
rect 9324 23866 9352 25094
rect 9600 24750 9628 25298
rect 9692 25294 9720 26182
rect 9772 25968 9824 25974
rect 9772 25910 9824 25916
rect 9956 25968 10008 25974
rect 9956 25910 10008 25916
rect 9680 25288 9732 25294
rect 9680 25230 9732 25236
rect 9680 24880 9732 24886
rect 9680 24822 9732 24828
rect 9588 24744 9640 24750
rect 9588 24686 9640 24692
rect 9312 23860 9364 23866
rect 9312 23802 9364 23808
rect 9600 23594 9628 24686
rect 9692 23662 9720 24822
rect 9784 24274 9812 25910
rect 9968 24818 9996 25910
rect 10152 24886 10180 26182
rect 10140 24880 10192 24886
rect 10140 24822 10192 24828
rect 9956 24812 10008 24818
rect 9956 24754 10008 24760
rect 9864 24676 9916 24682
rect 9864 24618 9916 24624
rect 9772 24268 9824 24274
rect 9772 24210 9824 24216
rect 9876 24206 9904 24618
rect 9864 24200 9916 24206
rect 9864 24142 9916 24148
rect 10244 23798 10272 36790
rect 10336 35290 10364 37810
rect 10428 37108 10456 38286
rect 12624 38276 12676 38282
rect 12624 38218 12676 38224
rect 12348 38208 12400 38214
rect 12348 38150 12400 38156
rect 10784 37868 10836 37874
rect 10784 37810 10836 37816
rect 11612 37868 11664 37874
rect 11612 37810 11664 37816
rect 10428 37080 10548 37108
rect 10416 36168 10468 36174
rect 10416 36110 10468 36116
rect 10324 35284 10376 35290
rect 10324 35226 10376 35232
rect 10324 35148 10376 35154
rect 10324 35090 10376 35096
rect 10336 32978 10364 35090
rect 10428 33998 10456 36110
rect 10416 33992 10468 33998
rect 10416 33934 10468 33940
rect 10520 33658 10548 37080
rect 10600 36712 10652 36718
rect 10600 36654 10652 36660
rect 10612 35154 10640 36654
rect 10692 36032 10744 36038
rect 10692 35974 10744 35980
rect 10704 35834 10732 35974
rect 10796 35834 10824 37810
rect 10968 37664 11020 37670
rect 10968 37606 11020 37612
rect 10876 37120 10928 37126
rect 10876 37062 10928 37068
rect 10888 36786 10916 37062
rect 10876 36780 10928 36786
rect 10876 36722 10928 36728
rect 10980 36106 11008 37606
rect 11244 36780 11296 36786
rect 11244 36722 11296 36728
rect 11256 36378 11284 36722
rect 11244 36372 11296 36378
rect 11244 36314 11296 36320
rect 10968 36100 11020 36106
rect 10968 36042 11020 36048
rect 10692 35828 10744 35834
rect 10692 35770 10744 35776
rect 10784 35828 10836 35834
rect 10784 35770 10836 35776
rect 10692 35624 10744 35630
rect 10692 35566 10744 35572
rect 10600 35148 10652 35154
rect 10600 35090 10652 35096
rect 10600 34944 10652 34950
rect 10600 34886 10652 34892
rect 10508 33652 10560 33658
rect 10508 33594 10560 33600
rect 10324 32972 10376 32978
rect 10324 32914 10376 32920
rect 10508 32224 10560 32230
rect 10508 32166 10560 32172
rect 10520 31754 10548 32166
rect 10508 31748 10560 31754
rect 10508 31690 10560 31696
rect 10508 26512 10560 26518
rect 10508 26454 10560 26460
rect 10520 25770 10548 26454
rect 10612 26234 10640 34886
rect 10704 34542 10732 35566
rect 10968 35148 11020 35154
rect 10968 35090 11020 35096
rect 10692 34536 10744 34542
rect 10692 34478 10744 34484
rect 10876 34468 10928 34474
rect 10876 34410 10928 34416
rect 10692 34400 10744 34406
rect 10692 34342 10744 34348
rect 10704 34066 10732 34342
rect 10692 34060 10744 34066
rect 10692 34002 10744 34008
rect 10888 31278 10916 34410
rect 10980 33454 11008 35090
rect 11256 35018 11284 36314
rect 11244 35012 11296 35018
rect 11244 34954 11296 34960
rect 11256 34610 11284 34954
rect 11244 34604 11296 34610
rect 11244 34546 11296 34552
rect 11152 34536 11204 34542
rect 11152 34478 11204 34484
rect 11164 33930 11192 34478
rect 11152 33924 11204 33930
rect 11152 33866 11204 33872
rect 10968 33448 11020 33454
rect 10968 33390 11020 33396
rect 11256 32910 11284 34546
rect 11244 32904 11296 32910
rect 11244 32846 11296 32852
rect 11060 32768 11112 32774
rect 11060 32710 11112 32716
rect 11520 32768 11572 32774
rect 11520 32710 11572 32716
rect 11072 32502 11100 32710
rect 11060 32496 11112 32502
rect 11060 32438 11112 32444
rect 10968 32428 11020 32434
rect 10968 32370 11020 32376
rect 10876 31272 10928 31278
rect 10876 31214 10928 31220
rect 10888 29714 10916 31214
rect 10980 30938 11008 32370
rect 11152 32224 11204 32230
rect 11152 32166 11204 32172
rect 11164 32026 11192 32166
rect 11060 32020 11112 32026
rect 11060 31962 11112 31968
rect 11152 32020 11204 32026
rect 11152 31962 11204 31968
rect 10968 30932 11020 30938
rect 10968 30874 11020 30880
rect 11072 29714 11100 31962
rect 11532 31958 11560 32710
rect 11520 31952 11572 31958
rect 11520 31894 11572 31900
rect 11532 31414 11560 31894
rect 11520 31408 11572 31414
rect 11520 31350 11572 31356
rect 11532 30802 11560 31350
rect 11520 30796 11572 30802
rect 11520 30738 11572 30744
rect 11152 30388 11204 30394
rect 11152 30330 11204 30336
rect 11164 30190 11192 30330
rect 11244 30252 11296 30258
rect 11244 30194 11296 30200
rect 11152 30184 11204 30190
rect 11152 30126 11204 30132
rect 11152 29776 11204 29782
rect 11256 29730 11284 30194
rect 11624 30054 11652 37810
rect 11980 37188 12032 37194
rect 11980 37130 12032 37136
rect 11992 36922 12020 37130
rect 12360 37126 12388 38150
rect 12256 37120 12308 37126
rect 12256 37062 12308 37068
rect 12348 37120 12400 37126
rect 12348 37062 12400 37068
rect 11980 36916 12032 36922
rect 11980 36858 12032 36864
rect 12072 36576 12124 36582
rect 12072 36518 12124 36524
rect 12084 36106 12112 36518
rect 12268 36310 12296 37062
rect 12636 36718 12664 38218
rect 13096 38010 13124 38286
rect 14096 38208 14148 38214
rect 14096 38150 14148 38156
rect 13084 38004 13136 38010
rect 13084 37946 13136 37952
rect 12808 37868 12860 37874
rect 12808 37810 12860 37816
rect 13452 37868 13504 37874
rect 13452 37810 13504 37816
rect 12624 36712 12676 36718
rect 12624 36654 12676 36660
rect 12256 36304 12308 36310
rect 12256 36246 12308 36252
rect 12072 36100 12124 36106
rect 12072 36042 12124 36048
rect 12164 35624 12216 35630
rect 12164 35566 12216 35572
rect 12176 35222 12204 35566
rect 12164 35216 12216 35222
rect 12164 35158 12216 35164
rect 12164 35080 12216 35086
rect 12164 35022 12216 35028
rect 11796 34944 11848 34950
rect 11796 34886 11848 34892
rect 11808 33590 11836 34886
rect 12072 34604 12124 34610
rect 12072 34546 12124 34552
rect 11980 34536 12032 34542
rect 11980 34478 12032 34484
rect 11992 33862 12020 34478
rect 11980 33856 12032 33862
rect 11980 33798 12032 33804
rect 11796 33584 11848 33590
rect 11796 33526 11848 33532
rect 12084 33114 12112 34546
rect 12176 34202 12204 35022
rect 12164 34196 12216 34202
rect 12164 34138 12216 34144
rect 12164 33856 12216 33862
rect 12164 33798 12216 33804
rect 12072 33108 12124 33114
rect 12072 33050 12124 33056
rect 12176 32842 12204 33798
rect 12268 33454 12296 36246
rect 12440 36236 12492 36242
rect 12440 36178 12492 36184
rect 12452 35170 12480 36178
rect 12452 35142 12572 35170
rect 12440 35080 12492 35086
rect 12440 35022 12492 35028
rect 12348 34944 12400 34950
rect 12348 34886 12400 34892
rect 12360 34678 12388 34886
rect 12348 34672 12400 34678
rect 12348 34614 12400 34620
rect 12256 33448 12308 33454
rect 12256 33390 12308 33396
rect 12164 32836 12216 32842
rect 12164 32778 12216 32784
rect 12072 32428 12124 32434
rect 12072 32370 12124 32376
rect 11704 32224 11756 32230
rect 11704 32166 11756 32172
rect 11716 31482 11744 32166
rect 11704 31476 11756 31482
rect 11704 31418 11756 31424
rect 11888 31340 11940 31346
rect 11888 31282 11940 31288
rect 11980 31340 12032 31346
rect 11980 31282 12032 31288
rect 11900 30938 11928 31282
rect 11888 30932 11940 30938
rect 11888 30874 11940 30880
rect 11992 30666 12020 31282
rect 11980 30660 12032 30666
rect 11980 30602 12032 30608
rect 11612 30048 11664 30054
rect 11612 29990 11664 29996
rect 11204 29724 11284 29730
rect 11152 29718 11284 29724
rect 10876 29708 10928 29714
rect 10876 29650 10928 29656
rect 11060 29708 11112 29714
rect 11164 29702 11284 29718
rect 11060 29650 11112 29656
rect 11152 29640 11204 29646
rect 11152 29582 11204 29588
rect 11164 29102 11192 29582
rect 11256 29306 11284 29702
rect 11244 29300 11296 29306
rect 11244 29242 11296 29248
rect 11704 29164 11756 29170
rect 11704 29106 11756 29112
rect 11152 29096 11204 29102
rect 11152 29038 11204 29044
rect 11244 28416 11296 28422
rect 11244 28358 11296 28364
rect 11336 28416 11388 28422
rect 11336 28358 11388 28364
rect 11256 28218 11284 28358
rect 11348 28218 11376 28358
rect 11244 28212 11296 28218
rect 11244 28154 11296 28160
rect 11336 28212 11388 28218
rect 11336 28154 11388 28160
rect 11060 27532 11112 27538
rect 11060 27474 11112 27480
rect 11072 26994 11100 27474
rect 11152 27328 11204 27334
rect 11152 27270 11204 27276
rect 11060 26988 11112 26994
rect 11060 26930 11112 26936
rect 11164 26382 11192 27270
rect 11256 27062 11284 28154
rect 11244 27056 11296 27062
rect 11244 26998 11296 27004
rect 11716 26994 11744 29106
rect 11796 29028 11848 29034
rect 11796 28970 11848 28976
rect 11808 27402 11836 28970
rect 11888 28416 11940 28422
rect 11888 28358 11940 28364
rect 11900 28082 11928 28358
rect 11888 28076 11940 28082
rect 11888 28018 11940 28024
rect 11796 27396 11848 27402
rect 11796 27338 11848 27344
rect 11704 26988 11756 26994
rect 11704 26930 11756 26936
rect 11796 26852 11848 26858
rect 11796 26794 11848 26800
rect 11428 26784 11480 26790
rect 11428 26726 11480 26732
rect 11244 26444 11296 26450
rect 11244 26386 11296 26392
rect 11152 26376 11204 26382
rect 11152 26318 11204 26324
rect 11256 26234 11284 26386
rect 11440 26314 11468 26726
rect 11808 26450 11836 26794
rect 11796 26444 11848 26450
rect 11796 26386 11848 26392
rect 11336 26308 11388 26314
rect 11336 26250 11388 26256
rect 11428 26308 11480 26314
rect 11428 26250 11480 26256
rect 10612 26206 10732 26234
rect 10508 25764 10560 25770
rect 10508 25706 10560 25712
rect 10520 25158 10548 25706
rect 10508 25152 10560 25158
rect 10508 25094 10560 25100
rect 10704 24954 10732 26206
rect 11164 26206 11284 26234
rect 10876 25900 10928 25906
rect 10876 25842 10928 25848
rect 10692 24948 10744 24954
rect 10692 24890 10744 24896
rect 10888 24682 10916 25842
rect 11164 25362 11192 26206
rect 11152 25356 11204 25362
rect 11152 25298 11204 25304
rect 10968 25288 11020 25294
rect 10968 25230 11020 25236
rect 10980 24682 11008 25230
rect 10876 24676 10928 24682
rect 10876 24618 10928 24624
rect 10968 24676 11020 24682
rect 10968 24618 11020 24624
rect 10784 24608 10836 24614
rect 10784 24550 10836 24556
rect 10796 23866 10824 24550
rect 10784 23860 10836 23866
rect 10784 23802 10836 23808
rect 10232 23792 10284 23798
rect 10232 23734 10284 23740
rect 9680 23656 9732 23662
rect 9680 23598 9732 23604
rect 9772 23656 9824 23662
rect 9772 23598 9824 23604
rect 9588 23588 9640 23594
rect 9588 23530 9640 23536
rect 9312 23520 9364 23526
rect 9312 23462 9364 23468
rect 9220 22976 9272 22982
rect 9220 22918 9272 22924
rect 9128 22636 9180 22642
rect 9128 22578 9180 22584
rect 8760 20868 8812 20874
rect 8760 20810 8812 20816
rect 8668 20800 8720 20806
rect 8668 20742 8720 20748
rect 8680 20602 8708 20742
rect 8668 20596 8720 20602
rect 8668 20538 8720 20544
rect 9140 20466 9168 22578
rect 9324 22030 9352 23462
rect 9600 23186 9628 23530
rect 9588 23180 9640 23186
rect 9588 23122 9640 23128
rect 9404 22568 9456 22574
rect 9404 22510 9456 22516
rect 9416 22234 9444 22510
rect 9404 22228 9456 22234
rect 9404 22170 9456 22176
rect 9312 22024 9364 22030
rect 9312 21966 9364 21972
rect 9496 22024 9548 22030
rect 9496 21966 9548 21972
rect 8484 20460 8536 20466
rect 8484 20402 8536 20408
rect 9128 20460 9180 20466
rect 9128 20402 9180 20408
rect 9508 19854 9536 21966
rect 9600 21078 9628 23122
rect 9692 22778 9720 23598
rect 9784 23254 9812 23598
rect 10600 23520 10652 23526
rect 10600 23462 10652 23468
rect 9772 23248 9824 23254
rect 9772 23190 9824 23196
rect 9680 22772 9732 22778
rect 9680 22714 9732 22720
rect 10048 22704 10100 22710
rect 10048 22646 10100 22652
rect 10060 22098 10088 22646
rect 10048 22092 10100 22098
rect 10048 22034 10100 22040
rect 10612 22030 10640 23462
rect 10784 23044 10836 23050
rect 10784 22986 10836 22992
rect 10796 22234 10824 22986
rect 10784 22228 10836 22234
rect 10784 22170 10836 22176
rect 10600 22024 10652 22030
rect 10600 21966 10652 21972
rect 10140 21548 10192 21554
rect 10140 21490 10192 21496
rect 9956 21344 10008 21350
rect 9956 21286 10008 21292
rect 9588 21072 9640 21078
rect 9588 21014 9640 21020
rect 9588 20936 9640 20942
rect 9588 20878 9640 20884
rect 8576 19848 8628 19854
rect 8576 19790 8628 19796
rect 9496 19848 9548 19854
rect 9496 19790 9548 19796
rect 8392 19712 8444 19718
rect 8392 19654 8444 19660
rect 8300 19440 8352 19446
rect 8300 19382 8352 19388
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 7012 18964 7064 18970
rect 7012 18906 7064 18912
rect 6000 18692 6052 18698
rect 6000 18634 6052 18640
rect 4874 18524 5182 18533
rect 4874 18522 4880 18524
rect 4936 18522 4960 18524
rect 5016 18522 5040 18524
rect 5096 18522 5120 18524
rect 5176 18522 5182 18524
rect 4936 18470 4938 18522
rect 5118 18470 5120 18522
rect 4874 18468 4880 18470
rect 4936 18468 4960 18470
rect 5016 18468 5040 18470
rect 5096 18468 5120 18470
rect 5176 18468 5182 18470
rect 4874 18459 5182 18468
rect 6012 18426 6040 18634
rect 6000 18420 6052 18426
rect 6000 18362 6052 18368
rect 6368 18284 6420 18290
rect 6368 18226 6420 18232
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 6092 17604 6144 17610
rect 6092 17546 6144 17552
rect 4874 17436 5182 17445
rect 4874 17434 4880 17436
rect 4936 17434 4960 17436
rect 5016 17434 5040 17436
rect 5096 17434 5120 17436
rect 5176 17434 5182 17436
rect 4936 17382 4938 17434
rect 5118 17382 5120 17434
rect 4874 17380 4880 17382
rect 4936 17380 4960 17382
rect 5016 17380 5040 17382
rect 5096 17380 5120 17382
rect 5176 17380 5182 17382
rect 4874 17371 5182 17380
rect 6104 17202 6132 17546
rect 5816 17196 5868 17202
rect 5816 17138 5868 17144
rect 6092 17196 6144 17202
rect 6092 17138 6144 17144
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4874 16348 5182 16357
rect 4874 16346 4880 16348
rect 4936 16346 4960 16348
rect 5016 16346 5040 16348
rect 5096 16346 5120 16348
rect 5176 16346 5182 16348
rect 4936 16294 4938 16346
rect 5118 16294 5120 16346
rect 4874 16292 4880 16294
rect 4936 16292 4960 16294
rect 5016 16292 5040 16294
rect 5096 16292 5120 16294
rect 5176 16292 5182 16294
rect 4874 16283 5182 16292
rect 5540 15904 5592 15910
rect 5540 15846 5592 15852
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4874 15260 5182 15269
rect 4874 15258 4880 15260
rect 4936 15258 4960 15260
rect 5016 15258 5040 15260
rect 5096 15258 5120 15260
rect 5176 15258 5182 15260
rect 4936 15206 4938 15258
rect 5118 15206 5120 15258
rect 4874 15204 4880 15206
rect 4936 15204 4960 15206
rect 5016 15204 5040 15206
rect 5096 15204 5120 15206
rect 5176 15204 5182 15206
rect 4874 15195 5182 15204
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 5552 14414 5580 15846
rect 5828 15502 5856 17138
rect 6092 16720 6144 16726
rect 6092 16662 6144 16668
rect 5816 15496 5868 15502
rect 5816 15438 5868 15444
rect 5540 14408 5592 14414
rect 5540 14350 5592 14356
rect 4874 14172 5182 14181
rect 4874 14170 4880 14172
rect 4936 14170 4960 14172
rect 5016 14170 5040 14172
rect 5096 14170 5120 14172
rect 5176 14170 5182 14172
rect 4936 14118 4938 14170
rect 5118 14118 5120 14170
rect 4874 14116 4880 14118
rect 4936 14116 4960 14118
rect 5016 14116 5040 14118
rect 5096 14116 5120 14118
rect 5176 14116 5182 14118
rect 4874 14107 5182 14116
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 2228 13456 2280 13462
rect 2228 13398 2280 13404
rect 5828 13326 5856 15438
rect 6104 14482 6132 16662
rect 6380 16454 6408 18226
rect 6644 17604 6696 17610
rect 6644 17546 6696 17552
rect 6552 17128 6604 17134
rect 6552 17070 6604 17076
rect 6368 16448 6420 16454
rect 6368 16390 6420 16396
rect 6564 15570 6592 17070
rect 6656 16522 6684 17546
rect 6736 17536 6788 17542
rect 6736 17478 6788 17484
rect 6920 17536 6972 17542
rect 6920 17478 6972 17484
rect 6748 17218 6776 17478
rect 6748 17190 6868 17218
rect 6840 17134 6868 17190
rect 6828 17128 6880 17134
rect 6828 17070 6880 17076
rect 6828 16992 6880 16998
rect 6932 16946 6960 17478
rect 6880 16940 6960 16946
rect 6828 16934 6960 16940
rect 6840 16918 6960 16934
rect 6840 16658 6868 16918
rect 6828 16652 6880 16658
rect 6828 16594 6880 16600
rect 7024 16590 7052 18906
rect 8312 18834 8340 19382
rect 8404 19310 8432 19654
rect 8588 19514 8616 19790
rect 9312 19712 9364 19718
rect 9312 19654 9364 19660
rect 8576 19508 8628 19514
rect 8576 19450 8628 19456
rect 9324 19446 9352 19654
rect 9312 19440 9364 19446
rect 9312 19382 9364 19388
rect 8392 19304 8444 19310
rect 8392 19246 8444 19252
rect 8300 18828 8352 18834
rect 8300 18770 8352 18776
rect 9404 18828 9456 18834
rect 9404 18770 9456 18776
rect 7288 18692 7340 18698
rect 7288 18634 7340 18640
rect 8392 18692 8444 18698
rect 8392 18634 8444 18640
rect 7300 18426 7328 18634
rect 7288 18420 7340 18426
rect 7288 18362 7340 18368
rect 7288 18284 7340 18290
rect 7288 18226 7340 18232
rect 7104 17740 7156 17746
rect 7104 17682 7156 17688
rect 7116 16794 7144 17682
rect 7104 16788 7156 16794
rect 7104 16730 7156 16736
rect 7012 16584 7064 16590
rect 7012 16526 7064 16532
rect 6644 16516 6696 16522
rect 6644 16458 6696 16464
rect 6920 16244 6972 16250
rect 6920 16186 6972 16192
rect 6552 15564 6604 15570
rect 6552 15506 6604 15512
rect 6552 15428 6604 15434
rect 6552 15370 6604 15376
rect 6564 15162 6592 15370
rect 6552 15156 6604 15162
rect 6552 15098 6604 15104
rect 6932 14618 6960 16186
rect 7116 15178 7144 16730
rect 7196 16652 7248 16658
rect 7196 16594 7248 16600
rect 7208 16046 7236 16594
rect 7196 16040 7248 16046
rect 7196 15982 7248 15988
rect 7116 15150 7236 15178
rect 7012 15020 7064 15026
rect 7012 14962 7064 14968
rect 6920 14612 6972 14618
rect 6920 14554 6972 14560
rect 6092 14476 6144 14482
rect 6092 14418 6144 14424
rect 5816 13320 5868 13326
rect 5816 13262 5868 13268
rect 4874 13084 5182 13093
rect 4874 13082 4880 13084
rect 4936 13082 4960 13084
rect 5016 13082 5040 13084
rect 5096 13082 5120 13084
rect 5176 13082 5182 13084
rect 4936 13030 4938 13082
rect 5118 13030 5120 13082
rect 4874 13028 4880 13030
rect 4936 13028 4960 13030
rect 5016 13028 5040 13030
rect 5096 13028 5120 13030
rect 5176 13028 5182 13030
rect 4874 13019 5182 13028
rect 6104 12850 6132 14418
rect 7024 14074 7052 14962
rect 7208 14958 7236 15150
rect 7196 14952 7248 14958
rect 7196 14894 7248 14900
rect 7012 14068 7064 14074
rect 7012 14010 7064 14016
rect 7012 13932 7064 13938
rect 7012 13874 7064 13880
rect 6092 12844 6144 12850
rect 6092 12786 6144 12792
rect 6552 12844 6604 12850
rect 6552 12786 6604 12792
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 6564 12306 6592 12786
rect 6828 12776 6880 12782
rect 6828 12718 6880 12724
rect 6840 12442 6868 12718
rect 7024 12646 7052 13874
rect 7104 13184 7156 13190
rect 7104 13126 7156 13132
rect 7116 12918 7144 13126
rect 7104 12912 7156 12918
rect 7104 12854 7156 12860
rect 7012 12640 7064 12646
rect 7012 12582 7064 12588
rect 6828 12436 6880 12442
rect 6828 12378 6880 12384
rect 6552 12300 6604 12306
rect 6552 12242 6604 12248
rect 6184 12232 6236 12238
rect 6184 12174 6236 12180
rect 4874 11996 5182 12005
rect 4874 11994 4880 11996
rect 4936 11994 4960 11996
rect 5016 11994 5040 11996
rect 5096 11994 5120 11996
rect 5176 11994 5182 11996
rect 4936 11942 4938 11994
rect 5118 11942 5120 11994
rect 4874 11940 4880 11942
rect 4936 11940 4960 11942
rect 5016 11940 5040 11942
rect 5096 11940 5120 11942
rect 5176 11940 5182 11942
rect 4874 11931 5182 11940
rect 6196 11898 6224 12174
rect 6184 11892 6236 11898
rect 6184 11834 6236 11840
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 6368 11008 6420 11014
rect 6368 10950 6420 10956
rect 4874 10908 5182 10917
rect 4874 10906 4880 10908
rect 4936 10906 4960 10908
rect 5016 10906 5040 10908
rect 5096 10906 5120 10908
rect 5176 10906 5182 10908
rect 4936 10854 4938 10906
rect 5118 10854 5120 10906
rect 4874 10852 4880 10854
rect 4936 10852 4960 10854
rect 5016 10852 5040 10854
rect 5096 10852 5120 10854
rect 5176 10852 5182 10854
rect 4874 10843 5182 10852
rect 1860 10804 1912 10810
rect 1860 10746 1912 10752
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 6380 9994 6408 10950
rect 6564 10742 6592 12242
rect 6920 11756 6972 11762
rect 6920 11698 6972 11704
rect 6644 11144 6696 11150
rect 6644 11086 6696 11092
rect 6552 10736 6604 10742
rect 6552 10678 6604 10684
rect 6564 10146 6592 10678
rect 6656 10538 6684 11086
rect 6644 10532 6696 10538
rect 6644 10474 6696 10480
rect 6472 10130 6592 10146
rect 6460 10124 6592 10130
rect 6512 10118 6592 10124
rect 6460 10066 6512 10072
rect 6368 9988 6420 9994
rect 6368 9930 6420 9936
rect 4874 9820 5182 9829
rect 4874 9818 4880 9820
rect 4936 9818 4960 9820
rect 5016 9818 5040 9820
rect 5096 9818 5120 9820
rect 5176 9818 5182 9820
rect 4936 9766 4938 9818
rect 5118 9766 5120 9818
rect 4874 9764 4880 9766
rect 4936 9764 4960 9766
rect 5016 9764 5040 9766
rect 5096 9764 5120 9766
rect 5176 9764 5182 9766
rect 4874 9755 5182 9764
rect 6932 9450 6960 11698
rect 7024 11694 7052 12582
rect 7104 12164 7156 12170
rect 7104 12106 7156 12112
rect 7012 11688 7064 11694
rect 7012 11630 7064 11636
rect 7024 10606 7052 11630
rect 7116 11354 7144 12106
rect 7208 11694 7236 14894
rect 7300 13326 7328 18226
rect 8404 17882 8432 18634
rect 9416 18290 9444 18770
rect 9220 18284 9272 18290
rect 9220 18226 9272 18232
rect 9404 18284 9456 18290
rect 9404 18226 9456 18232
rect 8392 17876 8444 17882
rect 8392 17818 8444 17824
rect 8760 17672 8812 17678
rect 8760 17614 8812 17620
rect 8772 17338 8800 17614
rect 9232 17542 9260 18226
rect 9508 17678 9536 19790
rect 9600 19786 9628 20878
rect 9968 20534 9996 21286
rect 9956 20528 10008 20534
rect 9956 20470 10008 20476
rect 10152 20058 10180 21490
rect 10888 21010 10916 24618
rect 11164 24274 11192 25298
rect 11348 24818 11376 26250
rect 11336 24812 11388 24818
rect 11336 24754 11388 24760
rect 11348 24342 11376 24754
rect 11336 24336 11388 24342
rect 11336 24278 11388 24284
rect 11152 24268 11204 24274
rect 11152 24210 11204 24216
rect 11704 24268 11756 24274
rect 11704 24210 11756 24216
rect 11336 24200 11388 24206
rect 11336 24142 11388 24148
rect 11348 23322 11376 24142
rect 11336 23316 11388 23322
rect 11336 23258 11388 23264
rect 11716 23202 11744 24210
rect 11992 24138 12020 30602
rect 12084 30258 12112 32370
rect 12164 32360 12216 32366
rect 12164 32302 12216 32308
rect 12176 30734 12204 32302
rect 12268 31890 12296 33390
rect 12452 32910 12480 35022
rect 12544 34066 12572 35142
rect 12636 35086 12664 36654
rect 12624 35080 12676 35086
rect 12624 35022 12676 35028
rect 12532 34060 12584 34066
rect 12532 34002 12584 34008
rect 12348 32904 12400 32910
rect 12348 32846 12400 32852
rect 12440 32904 12492 32910
rect 12440 32846 12492 32852
rect 12360 32434 12388 32846
rect 12348 32428 12400 32434
rect 12348 32370 12400 32376
rect 12348 32292 12400 32298
rect 12348 32234 12400 32240
rect 12360 32026 12388 32234
rect 12348 32020 12400 32026
rect 12348 31962 12400 31968
rect 12256 31884 12308 31890
rect 12256 31826 12308 31832
rect 12268 31278 12296 31826
rect 12452 31770 12480 32846
rect 12360 31742 12480 31770
rect 12256 31272 12308 31278
rect 12256 31214 12308 31220
rect 12360 31090 12388 31742
rect 12268 31062 12388 31090
rect 12164 30728 12216 30734
rect 12164 30670 12216 30676
rect 12072 30252 12124 30258
rect 12072 30194 12124 30200
rect 12268 30190 12296 31062
rect 12544 30802 12572 34002
rect 12624 33040 12676 33046
rect 12624 32982 12676 32988
rect 12636 32366 12664 32982
rect 12624 32360 12676 32366
rect 12624 32302 12676 32308
rect 12636 30870 12664 32302
rect 12624 30864 12676 30870
rect 12624 30806 12676 30812
rect 12532 30796 12584 30802
rect 12532 30738 12584 30744
rect 12544 30394 12572 30738
rect 12532 30388 12584 30394
rect 12532 30330 12584 30336
rect 12256 30184 12308 30190
rect 12440 30184 12492 30190
rect 12256 30126 12308 30132
rect 12360 30132 12440 30138
rect 12360 30126 12492 30132
rect 12360 30110 12480 30126
rect 12360 27538 12388 30110
rect 12544 28626 12572 30330
rect 12636 29186 12664 30806
rect 12636 29158 12756 29186
rect 12624 29096 12676 29102
rect 12624 29038 12676 29044
rect 12636 28762 12664 29038
rect 12624 28756 12676 28762
rect 12624 28698 12676 28704
rect 12532 28620 12584 28626
rect 12532 28562 12584 28568
rect 12544 27538 12572 28562
rect 12728 28014 12756 29158
rect 12716 28008 12768 28014
rect 12716 27950 12768 27956
rect 12164 27532 12216 27538
rect 12164 27474 12216 27480
rect 12348 27532 12400 27538
rect 12348 27474 12400 27480
rect 12532 27532 12584 27538
rect 12532 27474 12584 27480
rect 12176 27130 12204 27474
rect 12348 27396 12400 27402
rect 12348 27338 12400 27344
rect 12164 27124 12216 27130
rect 12164 27066 12216 27072
rect 12360 27062 12388 27338
rect 12348 27056 12400 27062
rect 12348 26998 12400 27004
rect 12544 26790 12572 27474
rect 12728 26926 12756 27950
rect 12716 26920 12768 26926
rect 12716 26862 12768 26868
rect 12532 26784 12584 26790
rect 12532 26726 12584 26732
rect 12820 26042 12848 37810
rect 13464 37466 13492 37810
rect 13452 37460 13504 37466
rect 13452 37402 13504 37408
rect 13464 36922 13492 37402
rect 13820 37324 13872 37330
rect 13820 37266 13872 37272
rect 13452 36916 13504 36922
rect 13452 36858 13504 36864
rect 13084 36712 13136 36718
rect 13084 36654 13136 36660
rect 13096 36174 13124 36654
rect 13464 36242 13492 36858
rect 13832 36854 13860 37266
rect 14108 36854 14136 38150
rect 14280 37868 14332 37874
rect 14280 37810 14332 37816
rect 13820 36848 13872 36854
rect 13820 36790 13872 36796
rect 14096 36848 14148 36854
rect 14096 36790 14148 36796
rect 13820 36712 13872 36718
rect 13820 36654 13872 36660
rect 13832 36310 13860 36654
rect 13820 36304 13872 36310
rect 13820 36246 13872 36252
rect 13452 36236 13504 36242
rect 13452 36178 13504 36184
rect 13084 36168 13136 36174
rect 13084 36110 13136 36116
rect 12992 36032 13044 36038
rect 12992 35974 13044 35980
rect 13004 35834 13032 35974
rect 13096 35894 13124 36110
rect 13096 35866 13216 35894
rect 12992 35828 13044 35834
rect 12992 35770 13044 35776
rect 13188 35630 13216 35866
rect 13176 35624 13228 35630
rect 13176 35566 13228 35572
rect 12992 34944 13044 34950
rect 12992 34886 13044 34892
rect 12900 33856 12952 33862
rect 12900 33798 12952 33804
rect 12912 33454 12940 33798
rect 13004 33590 13032 34886
rect 13188 34746 13216 35566
rect 13544 35556 13596 35562
rect 13544 35498 13596 35504
rect 13556 35086 13584 35498
rect 13832 35154 13860 36246
rect 14292 35894 14320 37810
rect 14372 37800 14424 37806
rect 14372 37742 14424 37748
rect 14464 37800 14516 37806
rect 14464 37742 14516 37748
rect 14384 37262 14412 37742
rect 14372 37256 14424 37262
rect 14372 37198 14424 37204
rect 14476 35894 14504 37742
rect 14660 37466 14688 38286
rect 14740 37732 14792 37738
rect 14740 37674 14792 37680
rect 14752 37466 14780 37674
rect 14648 37460 14700 37466
rect 14648 37402 14700 37408
rect 14740 37460 14792 37466
rect 14740 37402 14792 37408
rect 14924 37256 14976 37262
rect 14924 37198 14976 37204
rect 14936 36922 14964 37198
rect 14924 36916 14976 36922
rect 14924 36858 14976 36864
rect 14936 36106 14964 36858
rect 14924 36100 14976 36106
rect 14924 36042 14976 36048
rect 14292 35866 14412 35894
rect 14476 35866 14688 35894
rect 14280 35692 14332 35698
rect 14280 35634 14332 35640
rect 13912 35624 13964 35630
rect 13912 35566 13964 35572
rect 13820 35148 13872 35154
rect 13820 35090 13872 35096
rect 13544 35080 13596 35086
rect 13544 35022 13596 35028
rect 13452 35012 13504 35018
rect 13452 34954 13504 34960
rect 13464 34746 13492 34954
rect 13176 34740 13228 34746
rect 13176 34682 13228 34688
rect 13452 34740 13504 34746
rect 13452 34682 13504 34688
rect 13924 34542 13952 35566
rect 13912 34536 13964 34542
rect 13912 34478 13964 34484
rect 14188 34060 14240 34066
rect 14188 34002 14240 34008
rect 13912 33856 13964 33862
rect 13912 33798 13964 33804
rect 12992 33584 13044 33590
rect 12992 33526 13044 33532
rect 12900 33448 12952 33454
rect 12900 33390 12952 33396
rect 12912 32978 12940 33390
rect 12900 32972 12952 32978
rect 12900 32914 12952 32920
rect 13360 32768 13412 32774
rect 13360 32710 13412 32716
rect 13372 31822 13400 32710
rect 13360 31816 13412 31822
rect 13360 31758 13412 31764
rect 13820 31272 13872 31278
rect 13820 31214 13872 31220
rect 13636 30660 13688 30666
rect 13636 30602 13688 30608
rect 12900 30320 12952 30326
rect 12900 30262 12952 30268
rect 12912 29850 12940 30262
rect 12992 30252 13044 30258
rect 12992 30194 13044 30200
rect 12900 29844 12952 29850
rect 12900 29786 12952 29792
rect 13004 26194 13032 30194
rect 13648 29782 13676 30602
rect 13636 29776 13688 29782
rect 13636 29718 13688 29724
rect 13636 29504 13688 29510
rect 13636 29446 13688 29452
rect 13648 29238 13676 29446
rect 13636 29232 13688 29238
rect 13636 29174 13688 29180
rect 13832 29034 13860 31214
rect 13820 29028 13872 29034
rect 13820 28970 13872 28976
rect 13544 28416 13596 28422
rect 13544 28358 13596 28364
rect 13084 28076 13136 28082
rect 13084 28018 13136 28024
rect 13096 27334 13124 28018
rect 13084 27328 13136 27334
rect 13084 27270 13136 27276
rect 13096 26450 13124 27270
rect 13556 27062 13584 28358
rect 13728 28076 13780 28082
rect 13728 28018 13780 28024
rect 13636 27872 13688 27878
rect 13636 27814 13688 27820
rect 13648 27062 13676 27814
rect 13740 27402 13768 28018
rect 13728 27396 13780 27402
rect 13728 27338 13780 27344
rect 13740 27130 13768 27338
rect 13728 27124 13780 27130
rect 13728 27066 13780 27072
rect 13544 27056 13596 27062
rect 13544 26998 13596 27004
rect 13636 27056 13688 27062
rect 13636 26998 13688 27004
rect 13084 26444 13136 26450
rect 13084 26386 13136 26392
rect 12912 26166 13032 26194
rect 13820 26240 13872 26246
rect 13820 26182 13872 26188
rect 12808 26036 12860 26042
rect 12808 25978 12860 25984
rect 12164 25696 12216 25702
rect 12164 25638 12216 25644
rect 12072 25492 12124 25498
rect 12072 25434 12124 25440
rect 12084 24954 12112 25434
rect 12176 25226 12204 25638
rect 12164 25220 12216 25226
rect 12164 25162 12216 25168
rect 12072 24948 12124 24954
rect 12072 24890 12124 24896
rect 12164 24744 12216 24750
rect 12164 24686 12216 24692
rect 11980 24132 12032 24138
rect 11980 24074 12032 24080
rect 11888 24064 11940 24070
rect 11888 24006 11940 24012
rect 11796 23656 11848 23662
rect 11796 23598 11848 23604
rect 11532 23186 11744 23202
rect 11808 23186 11836 23598
rect 11520 23180 11744 23186
rect 11572 23174 11744 23180
rect 11520 23122 11572 23128
rect 11716 22642 11744 23174
rect 11796 23180 11848 23186
rect 11796 23122 11848 23128
rect 11900 22710 11928 24006
rect 11888 22704 11940 22710
rect 11888 22646 11940 22652
rect 11704 22636 11756 22642
rect 11704 22578 11756 22584
rect 11716 22166 11744 22578
rect 11704 22160 11756 22166
rect 11704 22102 11756 22108
rect 10876 21004 10928 21010
rect 10876 20946 10928 20952
rect 10784 20800 10836 20806
rect 10784 20742 10836 20748
rect 11612 20800 11664 20806
rect 11612 20742 11664 20748
rect 10796 20466 10824 20742
rect 11520 20596 11572 20602
rect 11520 20538 11572 20544
rect 10784 20460 10836 20466
rect 10784 20402 10836 20408
rect 10692 20392 10744 20398
rect 10692 20334 10744 20340
rect 10140 20052 10192 20058
rect 10140 19994 10192 20000
rect 9588 19780 9640 19786
rect 9588 19722 9640 19728
rect 9600 19378 9628 19722
rect 10600 19712 10652 19718
rect 10600 19654 10652 19660
rect 10612 19514 10640 19654
rect 10600 19508 10652 19514
rect 10600 19450 10652 19456
rect 9588 19372 9640 19378
rect 9588 19314 9640 19320
rect 10704 19242 10732 20334
rect 11532 19922 11560 20538
rect 11624 20534 11652 20742
rect 11612 20528 11664 20534
rect 11612 20470 11664 20476
rect 11716 20466 11744 22102
rect 11992 21078 12020 24074
rect 12176 23866 12204 24686
rect 12348 24268 12400 24274
rect 12348 24210 12400 24216
rect 12164 23860 12216 23866
rect 12164 23802 12216 23808
rect 12176 23254 12204 23802
rect 12360 23730 12388 24210
rect 12348 23724 12400 23730
rect 12348 23666 12400 23672
rect 12348 23588 12400 23594
rect 12348 23530 12400 23536
rect 12360 23474 12388 23530
rect 12532 23520 12584 23526
rect 12360 23446 12480 23474
rect 12532 23462 12584 23468
rect 12452 23254 12480 23446
rect 12164 23248 12216 23254
rect 12164 23190 12216 23196
rect 12440 23248 12492 23254
rect 12440 23190 12492 23196
rect 12544 23118 12572 23462
rect 12532 23112 12584 23118
rect 12532 23054 12584 23060
rect 12072 23044 12124 23050
rect 12072 22986 12124 22992
rect 12624 23044 12676 23050
rect 12624 22986 12676 22992
rect 12084 21690 12112 22986
rect 12440 22704 12492 22710
rect 12440 22646 12492 22652
rect 12452 22098 12480 22646
rect 12440 22092 12492 22098
rect 12440 22034 12492 22040
rect 12164 22024 12216 22030
rect 12164 21966 12216 21972
rect 12072 21684 12124 21690
rect 12072 21626 12124 21632
rect 12176 21554 12204 21966
rect 12440 21888 12492 21894
rect 12440 21830 12492 21836
rect 12164 21548 12216 21554
rect 12164 21490 12216 21496
rect 11980 21072 12032 21078
rect 11980 21014 12032 21020
rect 11704 20460 11756 20466
rect 11704 20402 11756 20408
rect 11060 19916 11112 19922
rect 11060 19858 11112 19864
rect 11520 19916 11572 19922
rect 11520 19858 11572 19864
rect 10692 19236 10744 19242
rect 10692 19178 10744 19184
rect 9864 18692 9916 18698
rect 9864 18634 9916 18640
rect 9680 18624 9732 18630
rect 9680 18566 9732 18572
rect 9496 17672 9548 17678
rect 9496 17614 9548 17620
rect 9220 17536 9272 17542
rect 9220 17478 9272 17484
rect 9692 17338 9720 18566
rect 9876 18426 9904 18634
rect 9864 18420 9916 18426
rect 9864 18362 9916 18368
rect 9772 18352 9824 18358
rect 9772 18294 9824 18300
rect 10140 18352 10192 18358
rect 10140 18294 10192 18300
rect 8208 17332 8260 17338
rect 8760 17332 8812 17338
rect 8260 17292 8524 17320
rect 8208 17274 8260 17280
rect 8208 16652 8260 16658
rect 8208 16594 8260 16600
rect 7932 16448 7984 16454
rect 7932 16390 7984 16396
rect 7840 16108 7892 16114
rect 7944 16096 7972 16390
rect 7892 16068 7972 16096
rect 7840 16050 7892 16056
rect 7944 15706 7972 16068
rect 7932 15700 7984 15706
rect 7932 15642 7984 15648
rect 7944 15162 7972 15642
rect 7932 15156 7984 15162
rect 7932 15098 7984 15104
rect 8116 15156 8168 15162
rect 8116 15098 8168 15104
rect 7472 14612 7524 14618
rect 7472 14554 7524 14560
rect 7380 14340 7432 14346
rect 7380 14282 7432 14288
rect 7392 13530 7420 14282
rect 7484 14074 7512 14554
rect 7472 14068 7524 14074
rect 7472 14010 7524 14016
rect 7380 13524 7432 13530
rect 7380 13466 7432 13472
rect 7288 13320 7340 13326
rect 7288 13262 7340 13268
rect 7300 11762 7328 13262
rect 7840 12164 7892 12170
rect 7840 12106 7892 12112
rect 7852 11898 7880 12106
rect 7840 11892 7892 11898
rect 7840 11834 7892 11840
rect 7288 11756 7340 11762
rect 7288 11698 7340 11704
rect 7932 11756 7984 11762
rect 7932 11698 7984 11704
rect 7196 11688 7248 11694
rect 7196 11630 7248 11636
rect 7104 11348 7156 11354
rect 7104 11290 7156 11296
rect 7012 10600 7064 10606
rect 7012 10542 7064 10548
rect 7104 9580 7156 9586
rect 7104 9522 7156 9528
rect 6920 9444 6972 9450
rect 6920 9386 6972 9392
rect 1584 9376 1636 9382
rect 1582 9344 1584 9353
rect 1636 9344 1638 9353
rect 1582 9279 1638 9288
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 7116 8838 7144 9522
rect 7208 9042 7236 11630
rect 7944 10674 7972 11698
rect 7840 10668 7892 10674
rect 7840 10610 7892 10616
rect 7932 10668 7984 10674
rect 7932 10610 7984 10616
rect 7656 10464 7708 10470
rect 7656 10406 7708 10412
rect 7668 9994 7696 10406
rect 7656 9988 7708 9994
rect 7656 9930 7708 9936
rect 7852 9926 7880 10610
rect 7840 9920 7892 9926
rect 7840 9862 7892 9868
rect 7852 9586 7880 9862
rect 7840 9580 7892 9586
rect 7840 9522 7892 9528
rect 7656 9512 7708 9518
rect 7656 9454 7708 9460
rect 7668 9042 7696 9454
rect 7196 9036 7248 9042
rect 7196 8978 7248 8984
rect 7656 9036 7708 9042
rect 7656 8978 7708 8984
rect 6092 8832 6144 8838
rect 6092 8774 6144 8780
rect 7104 8832 7156 8838
rect 7104 8774 7156 8780
rect 7380 8832 7432 8838
rect 7380 8774 7432 8780
rect 4874 8732 5182 8741
rect 4874 8730 4880 8732
rect 4936 8730 4960 8732
rect 5016 8730 5040 8732
rect 5096 8730 5120 8732
rect 5176 8730 5182 8732
rect 4936 8678 4938 8730
rect 5118 8678 5120 8730
rect 4874 8676 4880 8678
rect 4936 8676 4960 8678
rect 5016 8676 5040 8678
rect 5096 8676 5120 8678
rect 5176 8676 5182 8678
rect 4874 8667 5182 8676
rect 6104 8566 6132 8774
rect 6092 8560 6144 8566
rect 6092 8502 6144 8508
rect 5816 8492 5868 8498
rect 5816 8434 5868 8440
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 5828 8090 5856 8434
rect 7012 8356 7064 8362
rect 7012 8298 7064 8304
rect 5816 8084 5868 8090
rect 5816 8026 5868 8032
rect 7024 7818 7052 8298
rect 7116 7954 7144 8774
rect 7104 7948 7156 7954
rect 7104 7890 7156 7896
rect 7012 7812 7064 7818
rect 7012 7754 7064 7760
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 4874 7579 5182 7588
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 7024 5710 7052 7754
rect 7116 7546 7144 7890
rect 7392 7886 7420 8774
rect 7380 7880 7432 7886
rect 7380 7822 7432 7828
rect 7104 7540 7156 7546
rect 7104 7482 7156 7488
rect 7012 5704 7064 5710
rect 1582 5672 1638 5681
rect 7012 5646 7064 5652
rect 1582 5607 1638 5616
rect 1596 5574 1624 5607
rect 1584 5568 1636 5574
rect 1584 5510 1636 5516
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 7852 3058 7880 9522
rect 7944 9178 7972 10610
rect 7932 9172 7984 9178
rect 7932 9114 7984 9120
rect 7944 8974 7972 9114
rect 8128 9110 8156 15098
rect 8220 13734 8248 16594
rect 8300 15564 8352 15570
rect 8300 15506 8352 15512
rect 8312 14074 8340 15506
rect 8496 15502 8524 17292
rect 8760 17274 8812 17280
rect 9680 17332 9732 17338
rect 9680 17274 9732 17280
rect 9220 17128 9272 17134
rect 9220 17070 9272 17076
rect 9036 17060 9088 17066
rect 9036 17002 9088 17008
rect 9048 15910 9076 17002
rect 9232 16454 9260 17070
rect 9600 16794 9720 16810
rect 9588 16788 9720 16794
rect 9640 16782 9720 16788
rect 9588 16730 9640 16736
rect 9692 16574 9720 16782
rect 9600 16546 9720 16574
rect 9784 16574 9812 18294
rect 10152 17882 10180 18294
rect 10140 17876 10192 17882
rect 10140 17818 10192 17824
rect 10704 17746 10732 19178
rect 11072 18834 11100 19858
rect 12176 19854 12204 21490
rect 12452 20942 12480 21830
rect 12532 21072 12584 21078
rect 12532 21014 12584 21020
rect 12440 20936 12492 20942
rect 12440 20878 12492 20884
rect 12440 20528 12492 20534
rect 12440 20470 12492 20476
rect 12452 20058 12480 20470
rect 12440 20052 12492 20058
rect 12440 19994 12492 20000
rect 12164 19848 12216 19854
rect 12164 19790 12216 19796
rect 12440 19848 12492 19854
rect 12440 19790 12492 19796
rect 11612 19780 11664 19786
rect 11612 19722 11664 19728
rect 11624 18834 11652 19722
rect 11888 19372 11940 19378
rect 11888 19314 11940 19320
rect 11704 19168 11756 19174
rect 11704 19110 11756 19116
rect 11060 18828 11112 18834
rect 11060 18770 11112 18776
rect 11612 18828 11664 18834
rect 11612 18770 11664 18776
rect 11624 18426 11652 18770
rect 11152 18420 11204 18426
rect 11152 18362 11204 18368
rect 11612 18420 11664 18426
rect 11612 18362 11664 18368
rect 10692 17740 10744 17746
rect 10692 17682 10744 17688
rect 10508 17536 10560 17542
rect 10508 17478 10560 17484
rect 10520 17338 10548 17478
rect 10508 17332 10560 17338
rect 10508 17274 10560 17280
rect 10600 17128 10652 17134
rect 10600 17070 10652 17076
rect 9956 16992 10008 16998
rect 9956 16934 10008 16940
rect 9784 16546 9904 16574
rect 9404 16516 9456 16522
rect 9404 16458 9456 16464
rect 9220 16448 9272 16454
rect 9220 16390 9272 16396
rect 9232 16114 9260 16390
rect 9416 16250 9444 16458
rect 9404 16244 9456 16250
rect 9404 16186 9456 16192
rect 9220 16108 9272 16114
rect 9220 16050 9272 16056
rect 9600 16046 9628 16546
rect 9128 16040 9180 16046
rect 9128 15982 9180 15988
rect 9588 16040 9640 16046
rect 9588 15982 9640 15988
rect 9036 15904 9088 15910
rect 9036 15846 9088 15852
rect 8944 15564 8996 15570
rect 8944 15506 8996 15512
rect 8484 15496 8536 15502
rect 8484 15438 8536 15444
rect 8392 15360 8444 15366
rect 8392 15302 8444 15308
rect 8404 15026 8432 15302
rect 8956 15026 8984 15506
rect 9140 15162 9168 15982
rect 9404 15904 9456 15910
rect 9404 15846 9456 15852
rect 9416 15570 9444 15846
rect 9404 15564 9456 15570
rect 9404 15506 9456 15512
rect 9128 15156 9180 15162
rect 9128 15098 9180 15104
rect 8392 15020 8444 15026
rect 8392 14962 8444 14968
rect 8944 15020 8996 15026
rect 8944 14962 8996 14968
rect 8392 14408 8444 14414
rect 8392 14350 8444 14356
rect 8300 14068 8352 14074
rect 8300 14010 8352 14016
rect 8312 13938 8340 14010
rect 8300 13932 8352 13938
rect 8300 13874 8352 13880
rect 8208 13728 8260 13734
rect 8208 13670 8260 13676
rect 8404 13530 8432 14350
rect 8576 14272 8628 14278
rect 8576 14214 8628 14220
rect 9312 14272 9364 14278
rect 9312 14214 9364 14220
rect 8588 14006 8616 14214
rect 8576 14000 8628 14006
rect 8576 13942 8628 13948
rect 9036 14000 9088 14006
rect 9036 13942 9088 13948
rect 8392 13524 8444 13530
rect 8392 13466 8444 13472
rect 9048 13462 9076 13942
rect 8300 13456 8352 13462
rect 8300 13398 8352 13404
rect 9036 13456 9088 13462
rect 9036 13398 9088 13404
rect 8312 12918 8340 13398
rect 9324 13326 9352 14214
rect 8576 13320 8628 13326
rect 8576 13262 8628 13268
rect 9312 13320 9364 13326
rect 9312 13262 9364 13268
rect 8484 13252 8536 13258
rect 8484 13194 8536 13200
rect 8300 12912 8352 12918
rect 8300 12854 8352 12860
rect 8496 12782 8524 13194
rect 8484 12776 8536 12782
rect 8484 12718 8536 12724
rect 8496 12442 8524 12718
rect 8484 12436 8536 12442
rect 8484 12378 8536 12384
rect 8300 12368 8352 12374
rect 8300 12310 8352 12316
rect 8312 10606 8340 12310
rect 8588 12306 8616 13262
rect 9128 12640 9180 12646
rect 9128 12582 9180 12588
rect 8576 12300 8628 12306
rect 8576 12242 8628 12248
rect 8668 12096 8720 12102
rect 8668 12038 8720 12044
rect 8680 11150 8708 12038
rect 9140 11898 9168 12582
rect 9416 12374 9444 15506
rect 9876 15502 9904 16546
rect 9968 16182 9996 16934
rect 10140 16516 10192 16522
rect 10140 16458 10192 16464
rect 10152 16250 10180 16458
rect 10140 16244 10192 16250
rect 10140 16186 10192 16192
rect 9956 16176 10008 16182
rect 9956 16118 10008 16124
rect 9772 15496 9824 15502
rect 9772 15438 9824 15444
rect 9864 15496 9916 15502
rect 9864 15438 9916 15444
rect 9784 14958 9812 15438
rect 10048 15360 10100 15366
rect 10048 15302 10100 15308
rect 10324 15360 10376 15366
rect 10324 15302 10376 15308
rect 9772 14952 9824 14958
rect 9772 14894 9824 14900
rect 9784 14482 9812 14894
rect 9772 14476 9824 14482
rect 9772 14418 9824 14424
rect 9864 14476 9916 14482
rect 9864 14418 9916 14424
rect 9588 14068 9640 14074
rect 9588 14010 9640 14016
rect 9600 13870 9628 14010
rect 9588 13864 9640 13870
rect 9876 13818 9904 14418
rect 10060 14074 10088 15302
rect 10336 15026 10364 15302
rect 10324 15020 10376 15026
rect 10324 14962 10376 14968
rect 10612 14482 10640 17070
rect 10704 16794 10732 17682
rect 11164 17678 11192 18362
rect 11152 17672 11204 17678
rect 11152 17614 11204 17620
rect 11716 17610 11744 19110
rect 11900 18970 11928 19314
rect 11888 18964 11940 18970
rect 11888 18906 11940 18912
rect 12452 18834 12480 19790
rect 12440 18828 12492 18834
rect 12440 18770 12492 18776
rect 12164 18624 12216 18630
rect 12164 18566 12216 18572
rect 12072 18080 12124 18086
rect 12072 18022 12124 18028
rect 12084 17610 12112 18022
rect 12176 17882 12204 18566
rect 12164 17876 12216 17882
rect 12164 17818 12216 17824
rect 10784 17604 10836 17610
rect 10784 17546 10836 17552
rect 11704 17604 11756 17610
rect 11704 17546 11756 17552
rect 12072 17604 12124 17610
rect 12072 17546 12124 17552
rect 10692 16788 10744 16794
rect 10692 16730 10744 16736
rect 10796 16590 10824 17546
rect 12176 17338 12204 17818
rect 12164 17332 12216 17338
rect 12164 17274 12216 17280
rect 12440 17196 12492 17202
rect 12440 17138 12492 17144
rect 10784 16584 10836 16590
rect 10784 16526 10836 16532
rect 10796 16114 10824 16526
rect 11980 16448 12032 16454
rect 11980 16390 12032 16396
rect 12256 16448 12308 16454
rect 12256 16390 12308 16396
rect 10784 16108 10836 16114
rect 10784 16050 10836 16056
rect 11152 15904 11204 15910
rect 11152 15846 11204 15852
rect 11164 15706 11192 15846
rect 11152 15700 11204 15706
rect 11152 15642 11204 15648
rect 11992 15434 12020 16390
rect 12268 16250 12296 16390
rect 12256 16244 12308 16250
rect 12256 16186 12308 16192
rect 12452 16114 12480 17138
rect 12440 16108 12492 16114
rect 12440 16050 12492 16056
rect 11980 15428 12032 15434
rect 11980 15370 12032 15376
rect 11704 15020 11756 15026
rect 11704 14962 11756 14968
rect 11716 14618 11744 14962
rect 11888 14816 11940 14822
rect 11888 14758 11940 14764
rect 12256 14816 12308 14822
rect 12256 14758 12308 14764
rect 11704 14612 11756 14618
rect 11704 14554 11756 14560
rect 10968 14544 11020 14550
rect 10968 14486 11020 14492
rect 10600 14476 10652 14482
rect 10600 14418 10652 14424
rect 10692 14340 10744 14346
rect 10692 14282 10744 14288
rect 10704 14074 10732 14282
rect 10980 14278 11008 14486
rect 11244 14408 11296 14414
rect 11244 14350 11296 14356
rect 10784 14272 10836 14278
rect 10784 14214 10836 14220
rect 10968 14272 11020 14278
rect 10968 14214 11020 14220
rect 10048 14068 10100 14074
rect 10048 14010 10100 14016
rect 10692 14068 10744 14074
rect 10692 14010 10744 14016
rect 9640 13812 9720 13818
rect 9588 13806 9720 13812
rect 9600 13790 9720 13806
rect 9600 13741 9628 13790
rect 9692 13530 9720 13790
rect 9784 13790 9904 13818
rect 9784 13734 9812 13790
rect 9772 13728 9824 13734
rect 9772 13670 9824 13676
rect 9680 13524 9732 13530
rect 9680 13466 9732 13472
rect 9784 12782 9812 13670
rect 10060 13326 10088 14010
rect 10508 13932 10560 13938
rect 10508 13874 10560 13880
rect 10048 13320 10100 13326
rect 10048 13262 10100 13268
rect 10060 12986 10088 13262
rect 10520 12986 10548 13874
rect 10600 13728 10652 13734
rect 10600 13670 10652 13676
rect 10612 13394 10640 13670
rect 10600 13388 10652 13394
rect 10600 13330 10652 13336
rect 10600 13252 10652 13258
rect 10600 13194 10652 13200
rect 10048 12980 10100 12986
rect 10048 12922 10100 12928
rect 10508 12980 10560 12986
rect 10508 12922 10560 12928
rect 9496 12776 9548 12782
rect 9496 12718 9548 12724
rect 9772 12776 9824 12782
rect 9772 12718 9824 12724
rect 9404 12368 9456 12374
rect 9404 12310 9456 12316
rect 9508 12238 9536 12718
rect 9496 12232 9548 12238
rect 9496 12174 9548 12180
rect 9588 12232 9640 12238
rect 9588 12174 9640 12180
rect 9128 11892 9180 11898
rect 9128 11834 9180 11840
rect 9600 11830 9628 12174
rect 9680 12096 9732 12102
rect 9680 12038 9732 12044
rect 9692 11898 9720 12038
rect 9680 11892 9732 11898
rect 9680 11834 9732 11840
rect 9588 11824 9640 11830
rect 9588 11766 9640 11772
rect 8760 11552 8812 11558
rect 8760 11494 8812 11500
rect 8668 11144 8720 11150
rect 8668 11086 8720 11092
rect 8392 10804 8444 10810
rect 8392 10746 8444 10752
rect 8300 10600 8352 10606
rect 8300 10542 8352 10548
rect 8312 9586 8340 10542
rect 8404 10198 8432 10746
rect 8772 10742 8800 11494
rect 9600 11150 9628 11766
rect 9784 11218 9812 12718
rect 10612 12714 10640 13194
rect 10796 12986 10824 14214
rect 11060 14068 11112 14074
rect 11060 14010 11112 14016
rect 11072 12986 11100 14010
rect 10784 12980 10836 12986
rect 10784 12922 10836 12928
rect 11060 12980 11112 12986
rect 11060 12922 11112 12928
rect 11060 12844 11112 12850
rect 11060 12786 11112 12792
rect 10600 12708 10652 12714
rect 10600 12650 10652 12656
rect 10232 11892 10284 11898
rect 10232 11834 10284 11840
rect 9772 11212 9824 11218
rect 9772 11154 9824 11160
rect 9588 11144 9640 11150
rect 9588 11086 9640 11092
rect 9496 11008 9548 11014
rect 9496 10950 9548 10956
rect 9508 10742 9536 10950
rect 8760 10736 8812 10742
rect 8760 10678 8812 10684
rect 9496 10736 9548 10742
rect 9496 10678 9548 10684
rect 8392 10192 8444 10198
rect 8392 10134 8444 10140
rect 8392 10056 8444 10062
rect 8392 9998 8444 10004
rect 8404 9722 8432 9998
rect 8392 9716 8444 9722
rect 8392 9658 8444 9664
rect 8300 9580 8352 9586
rect 8300 9522 8352 9528
rect 8208 9512 8260 9518
rect 8208 9454 8260 9460
rect 8116 9104 8168 9110
rect 8116 9046 8168 9052
rect 8220 8974 8248 9454
rect 7932 8968 7984 8974
rect 7932 8910 7984 8916
rect 8208 8968 8260 8974
rect 8208 8910 8260 8916
rect 8024 8832 8076 8838
rect 8024 8774 8076 8780
rect 8036 7818 8064 8774
rect 8220 8634 8248 8910
rect 8208 8628 8260 8634
rect 8208 8570 8260 8576
rect 8312 7954 8340 9522
rect 9784 9450 9812 11154
rect 10140 11144 10192 11150
rect 10140 11086 10192 11092
rect 10152 10810 10180 11086
rect 10244 10810 10272 11834
rect 10612 11694 10640 12650
rect 11072 12374 11100 12786
rect 11256 12782 11284 14350
rect 11900 14006 11928 14758
rect 12268 14482 12296 14758
rect 12256 14476 12308 14482
rect 12256 14418 12308 14424
rect 12164 14340 12216 14346
rect 12164 14282 12216 14288
rect 12176 14074 12204 14282
rect 12164 14068 12216 14074
rect 12164 14010 12216 14016
rect 11888 14000 11940 14006
rect 11888 13942 11940 13948
rect 12176 13530 12204 14010
rect 12164 13524 12216 13530
rect 12164 13466 12216 13472
rect 12268 12850 12296 14418
rect 12440 13728 12492 13734
rect 12440 13670 12492 13676
rect 12544 13682 12572 21014
rect 12636 21010 12664 22986
rect 12820 21894 12848 25978
rect 12808 21888 12860 21894
rect 12808 21830 12860 21836
rect 12624 21004 12676 21010
rect 12624 20946 12676 20952
rect 12636 19530 12664 20946
rect 12912 20602 12940 26166
rect 13832 25906 13860 26182
rect 13820 25900 13872 25906
rect 13820 25842 13872 25848
rect 13728 25832 13780 25838
rect 13728 25774 13780 25780
rect 13740 25294 13768 25774
rect 13728 25288 13780 25294
rect 13728 25230 13780 25236
rect 12992 24744 13044 24750
rect 12992 24686 13044 24692
rect 13176 24744 13228 24750
rect 13176 24686 13228 24692
rect 13004 22001 13032 24686
rect 13084 23248 13136 23254
rect 13084 23190 13136 23196
rect 13096 22098 13124 23190
rect 13188 23186 13216 24686
rect 13544 24608 13596 24614
rect 13544 24550 13596 24556
rect 13556 24206 13584 24550
rect 13544 24200 13596 24206
rect 13544 24142 13596 24148
rect 13268 24064 13320 24070
rect 13268 24006 13320 24012
rect 13280 23798 13308 24006
rect 13268 23792 13320 23798
rect 13268 23734 13320 23740
rect 13924 23322 13952 33798
rect 14200 33318 14228 34002
rect 14188 33312 14240 33318
rect 14188 33254 14240 33260
rect 14200 32960 14228 33254
rect 14292 33114 14320 35634
rect 14280 33108 14332 33114
rect 14280 33050 14332 33056
rect 14200 32932 14320 32960
rect 14292 31890 14320 32932
rect 14280 31884 14332 31890
rect 14280 31826 14332 31832
rect 14004 31680 14056 31686
rect 14004 31622 14056 31628
rect 14016 23662 14044 31622
rect 14292 30190 14320 31826
rect 14280 30184 14332 30190
rect 14280 30126 14332 30132
rect 14096 28960 14148 28966
rect 14096 28902 14148 28908
rect 14108 28150 14136 28902
rect 14188 28552 14240 28558
rect 14188 28494 14240 28500
rect 14200 28218 14228 28494
rect 14188 28212 14240 28218
rect 14188 28154 14240 28160
rect 14096 28144 14148 28150
rect 14096 28086 14148 28092
rect 14188 27328 14240 27334
rect 14188 27270 14240 27276
rect 14200 25974 14228 27270
rect 14188 25968 14240 25974
rect 14188 25910 14240 25916
rect 14384 25158 14412 35866
rect 14464 35488 14516 35494
rect 14464 35430 14516 35436
rect 14476 32230 14504 35430
rect 14556 35148 14608 35154
rect 14556 35090 14608 35096
rect 14568 34678 14596 35090
rect 14556 34672 14608 34678
rect 14556 34614 14608 34620
rect 14660 34066 14688 35866
rect 14648 34060 14700 34066
rect 14648 34002 14700 34008
rect 14464 32224 14516 32230
rect 14464 32166 14516 32172
rect 15028 32026 15056 38286
rect 15200 38276 15252 38282
rect 15200 38218 15252 38224
rect 15108 37324 15160 37330
rect 15108 37266 15160 37272
rect 15120 36718 15148 37266
rect 15212 36786 15240 38218
rect 15764 38010 15792 38286
rect 18604 38276 18656 38282
rect 18604 38218 18656 38224
rect 17132 38208 17184 38214
rect 17132 38150 17184 38156
rect 18144 38208 18196 38214
rect 18144 38150 18196 38156
rect 15752 38004 15804 38010
rect 15752 37946 15804 37952
rect 17144 37942 17172 38150
rect 17132 37936 17184 37942
rect 17132 37878 17184 37884
rect 15292 37868 15344 37874
rect 15292 37810 15344 37816
rect 15200 36780 15252 36786
rect 15200 36722 15252 36728
rect 15108 36712 15160 36718
rect 15108 36654 15160 36660
rect 15108 35624 15160 35630
rect 15108 35566 15160 35572
rect 15120 33402 15148 35566
rect 15304 34202 15332 37810
rect 16856 37800 16908 37806
rect 16856 37742 16908 37748
rect 16028 37188 16080 37194
rect 16028 37130 16080 37136
rect 15384 37120 15436 37126
rect 15384 37062 15436 37068
rect 15396 35698 15424 37062
rect 16040 36922 16068 37130
rect 16868 37126 16896 37742
rect 17040 37188 17092 37194
rect 17040 37130 17092 37136
rect 16856 37120 16908 37126
rect 16856 37062 16908 37068
rect 16028 36916 16080 36922
rect 16028 36858 16080 36864
rect 17052 36378 17080 37130
rect 17316 37120 17368 37126
rect 17316 37062 17368 37068
rect 17960 37120 18012 37126
rect 17960 37062 18012 37068
rect 17132 36712 17184 36718
rect 17132 36654 17184 36660
rect 17040 36372 17092 36378
rect 17040 36314 17092 36320
rect 16028 36236 16080 36242
rect 16028 36178 16080 36184
rect 15568 36032 15620 36038
rect 15568 35974 15620 35980
rect 15580 35834 15608 35974
rect 15568 35828 15620 35834
rect 15568 35770 15620 35776
rect 15384 35692 15436 35698
rect 15384 35634 15436 35640
rect 15936 35692 15988 35698
rect 15936 35634 15988 35640
rect 15568 35012 15620 35018
rect 15568 34954 15620 34960
rect 15580 34746 15608 34954
rect 15948 34950 15976 35634
rect 15936 34944 15988 34950
rect 15936 34886 15988 34892
rect 15568 34740 15620 34746
rect 15568 34682 15620 34688
rect 15292 34196 15344 34202
rect 15292 34138 15344 34144
rect 15948 33998 15976 34886
rect 16040 34474 16068 36178
rect 17040 36168 17092 36174
rect 17040 36110 17092 36116
rect 16120 35488 16172 35494
rect 16120 35430 16172 35436
rect 16396 35488 16448 35494
rect 16396 35430 16448 35436
rect 16028 34468 16080 34474
rect 16028 34410 16080 34416
rect 16040 34066 16068 34410
rect 16132 34406 16160 35430
rect 16304 35012 16356 35018
rect 16304 34954 16356 34960
rect 16316 34746 16344 34954
rect 16304 34740 16356 34746
rect 16304 34682 16356 34688
rect 16408 34610 16436 35430
rect 16764 35148 16816 35154
rect 16764 35090 16816 35096
rect 16396 34604 16448 34610
rect 16396 34546 16448 34552
rect 16120 34400 16172 34406
rect 16120 34342 16172 34348
rect 16028 34060 16080 34066
rect 16028 34002 16080 34008
rect 15936 33992 15988 33998
rect 15936 33934 15988 33940
rect 15568 33856 15620 33862
rect 15568 33798 15620 33804
rect 15120 33374 15240 33402
rect 15108 33312 15160 33318
rect 15108 33254 15160 33260
rect 15120 33114 15148 33254
rect 15108 33108 15160 33114
rect 15108 33050 15160 33056
rect 15212 32978 15240 33374
rect 15580 33046 15608 33798
rect 16040 33538 16068 34002
rect 16580 33856 16632 33862
rect 16580 33798 16632 33804
rect 16592 33658 16620 33798
rect 16580 33652 16632 33658
rect 16580 33594 16632 33600
rect 16040 33510 16160 33538
rect 16028 33448 16080 33454
rect 16028 33390 16080 33396
rect 15568 33040 15620 33046
rect 15568 32982 15620 32988
rect 15200 32972 15252 32978
rect 15200 32914 15252 32920
rect 15212 32858 15240 32914
rect 15120 32830 15240 32858
rect 15016 32020 15068 32026
rect 15016 31962 15068 31968
rect 15120 30870 15148 32830
rect 16040 32774 16068 33390
rect 15200 32768 15252 32774
rect 15200 32710 15252 32716
rect 16028 32768 16080 32774
rect 16028 32710 16080 32716
rect 15212 32570 15240 32710
rect 15200 32564 15252 32570
rect 15200 32506 15252 32512
rect 15200 32360 15252 32366
rect 15252 32320 15332 32348
rect 15200 32302 15252 32308
rect 15304 31414 15332 32320
rect 16040 31822 16068 32710
rect 16132 31890 16160 33510
rect 16212 33448 16264 33454
rect 16212 33390 16264 33396
rect 16672 33448 16724 33454
rect 16776 33436 16804 35090
rect 17052 34134 17080 36110
rect 17040 34128 17092 34134
rect 17040 34070 17092 34076
rect 16856 33856 16908 33862
rect 16856 33798 16908 33804
rect 16724 33408 16804 33436
rect 16672 33390 16724 33396
rect 16120 31884 16172 31890
rect 16120 31826 16172 31832
rect 16028 31816 16080 31822
rect 16028 31758 16080 31764
rect 15568 31680 15620 31686
rect 15568 31622 15620 31628
rect 16028 31680 16080 31686
rect 16028 31622 16080 31628
rect 15292 31408 15344 31414
rect 15292 31350 15344 31356
rect 15108 30864 15160 30870
rect 15108 30806 15160 30812
rect 14832 30796 14884 30802
rect 14832 30738 14884 30744
rect 14844 30326 14872 30738
rect 15580 30734 15608 31622
rect 16040 31414 16068 31622
rect 16028 31408 16080 31414
rect 16028 31350 16080 31356
rect 16040 30938 16068 31350
rect 16132 30938 16160 31826
rect 16028 30932 16080 30938
rect 16028 30874 16080 30880
rect 16120 30932 16172 30938
rect 16120 30874 16172 30880
rect 15568 30728 15620 30734
rect 15568 30670 15620 30676
rect 14832 30320 14884 30326
rect 14832 30262 14884 30268
rect 15106 30288 15162 30297
rect 14924 30252 14976 30258
rect 15106 30223 15108 30232
rect 14924 30194 14976 30200
rect 15160 30223 15162 30232
rect 15752 30252 15804 30258
rect 15108 30194 15160 30200
rect 15752 30194 15804 30200
rect 14648 29572 14700 29578
rect 14648 29514 14700 29520
rect 14660 29306 14688 29514
rect 14648 29300 14700 29306
rect 14648 29242 14700 29248
rect 14556 29096 14608 29102
rect 14556 29038 14608 29044
rect 14568 27606 14596 29038
rect 14660 28558 14688 29242
rect 14648 28552 14700 28558
rect 14648 28494 14700 28500
rect 14832 28484 14884 28490
rect 14832 28426 14884 28432
rect 14648 28416 14700 28422
rect 14648 28358 14700 28364
rect 14740 28416 14792 28422
rect 14740 28358 14792 28364
rect 14660 28218 14688 28358
rect 14648 28212 14700 28218
rect 14648 28154 14700 28160
rect 14752 28150 14780 28358
rect 14740 28144 14792 28150
rect 14740 28086 14792 28092
rect 14556 27600 14608 27606
rect 14556 27542 14608 27548
rect 14556 27464 14608 27470
rect 14556 27406 14608 27412
rect 14568 27130 14596 27406
rect 14556 27124 14608 27130
rect 14556 27066 14608 27072
rect 14556 25696 14608 25702
rect 14556 25638 14608 25644
rect 14568 25362 14596 25638
rect 14556 25356 14608 25362
rect 14556 25298 14608 25304
rect 14648 25356 14700 25362
rect 14648 25298 14700 25304
rect 14660 25226 14688 25298
rect 14648 25220 14700 25226
rect 14648 25162 14700 25168
rect 14372 25152 14424 25158
rect 14372 25094 14424 25100
rect 14740 24880 14792 24886
rect 14740 24822 14792 24828
rect 14464 24676 14516 24682
rect 14464 24618 14516 24624
rect 14476 24206 14504 24618
rect 14464 24200 14516 24206
rect 14464 24142 14516 24148
rect 14372 24064 14424 24070
rect 14372 24006 14424 24012
rect 14384 23730 14412 24006
rect 14372 23724 14424 23730
rect 14372 23666 14424 23672
rect 14004 23656 14056 23662
rect 14004 23598 14056 23604
rect 13912 23316 13964 23322
rect 13912 23258 13964 23264
rect 13176 23180 13228 23186
rect 13228 23140 13308 23168
rect 13176 23122 13228 23128
rect 13280 22778 13308 23140
rect 13924 22982 13952 23258
rect 13912 22976 13964 22982
rect 13912 22918 13964 22924
rect 13268 22772 13320 22778
rect 13268 22714 13320 22720
rect 13084 22092 13136 22098
rect 13280 22094 13308 22714
rect 13912 22636 13964 22642
rect 13912 22578 13964 22584
rect 13084 22034 13136 22040
rect 13188 22066 13308 22094
rect 12990 21992 13046 22001
rect 12990 21927 13046 21936
rect 12992 21888 13044 21894
rect 12992 21830 13044 21836
rect 13004 21622 13032 21830
rect 12992 21616 13044 21622
rect 12992 21558 13044 21564
rect 12900 20596 12952 20602
rect 12900 20538 12952 20544
rect 13096 19922 13124 22034
rect 13188 22030 13216 22066
rect 13176 22024 13228 22030
rect 13176 21966 13228 21972
rect 13266 21992 13322 22001
rect 13266 21927 13322 21936
rect 13280 21486 13308 21927
rect 13924 21690 13952 22578
rect 14016 22506 14044 23598
rect 14004 22500 14056 22506
rect 14004 22442 14056 22448
rect 14096 22432 14148 22438
rect 14096 22374 14148 22380
rect 14108 22234 14136 22374
rect 14096 22228 14148 22234
rect 14096 22170 14148 22176
rect 14476 22094 14504 24142
rect 14752 23866 14780 24822
rect 14740 23860 14792 23866
rect 14740 23802 14792 23808
rect 14648 22704 14700 22710
rect 14648 22646 14700 22652
rect 14384 22066 14504 22094
rect 14096 22024 14148 22030
rect 14096 21966 14148 21972
rect 13912 21684 13964 21690
rect 13912 21626 13964 21632
rect 13268 21480 13320 21486
rect 13268 21422 13320 21428
rect 13452 21480 13504 21486
rect 13452 21422 13504 21428
rect 13464 20806 13492 21422
rect 13452 20800 13504 20806
rect 13452 20742 13504 20748
rect 13464 20602 13492 20742
rect 13452 20596 13504 20602
rect 13452 20538 13504 20544
rect 12808 19916 12860 19922
rect 12808 19858 12860 19864
rect 13084 19916 13136 19922
rect 13084 19858 13136 19864
rect 12636 19502 12756 19530
rect 12624 19440 12676 19446
rect 12624 19382 12676 19388
rect 12636 18222 12664 19382
rect 12728 19310 12756 19502
rect 12716 19304 12768 19310
rect 12716 19246 12768 19252
rect 12624 18216 12676 18222
rect 12624 18158 12676 18164
rect 12636 17746 12664 18158
rect 12624 17740 12676 17746
rect 12624 17682 12676 17688
rect 12820 17116 12848 19858
rect 13464 19854 13492 20538
rect 14108 20398 14136 21966
rect 14384 21554 14412 22066
rect 14372 21548 14424 21554
rect 14372 21490 14424 21496
rect 14384 20942 14412 21490
rect 14280 20936 14332 20942
rect 14280 20878 14332 20884
rect 14372 20936 14424 20942
rect 14372 20878 14424 20884
rect 14096 20392 14148 20398
rect 14096 20334 14148 20340
rect 13452 19848 13504 19854
rect 13452 19790 13504 19796
rect 13728 19712 13780 19718
rect 13728 19654 13780 19660
rect 13740 19514 13768 19654
rect 13728 19508 13780 19514
rect 13728 19450 13780 19456
rect 14108 19446 14136 20334
rect 14292 20058 14320 20878
rect 14280 20052 14332 20058
rect 14280 19994 14332 20000
rect 14096 19440 14148 19446
rect 14096 19382 14148 19388
rect 14384 19334 14412 20878
rect 14464 20800 14516 20806
rect 14464 20742 14516 20748
rect 14476 20534 14504 20742
rect 14464 20528 14516 20534
rect 14464 20470 14516 20476
rect 14464 19780 14516 19786
rect 14464 19722 14516 19728
rect 14476 19378 14504 19722
rect 13636 19304 13688 19310
rect 13636 19246 13688 19252
rect 13728 19304 13780 19310
rect 13728 19246 13780 19252
rect 14292 19306 14412 19334
rect 14464 19372 14516 19378
rect 14464 19314 14516 19320
rect 12900 19168 12952 19174
rect 12900 19110 12952 19116
rect 12912 18358 12940 19110
rect 13544 18760 13596 18766
rect 13544 18702 13596 18708
rect 13360 18692 13412 18698
rect 13360 18634 13412 18640
rect 12992 18624 13044 18630
rect 12992 18566 13044 18572
rect 13004 18358 13032 18566
rect 12900 18352 12952 18358
rect 12900 18294 12952 18300
rect 12992 18352 13044 18358
rect 12992 18294 13044 18300
rect 13372 17814 13400 18634
rect 13556 18426 13584 18702
rect 13544 18420 13596 18426
rect 13544 18362 13596 18368
rect 13360 17808 13412 17814
rect 13360 17750 13412 17756
rect 13372 17134 13400 17750
rect 13648 17746 13676 19246
rect 13740 18970 13768 19246
rect 13728 18964 13780 18970
rect 13728 18906 13780 18912
rect 13728 18828 13780 18834
rect 13728 18770 13780 18776
rect 13636 17740 13688 17746
rect 13636 17682 13688 17688
rect 13648 17338 13676 17682
rect 13636 17332 13688 17338
rect 13636 17274 13688 17280
rect 12900 17128 12952 17134
rect 12820 17088 12900 17116
rect 12900 17070 12952 17076
rect 13360 17128 13412 17134
rect 13648 17116 13676 17274
rect 13740 17218 13768 18770
rect 14292 18766 14320 19306
rect 14476 18766 14504 19314
rect 14280 18760 14332 18766
rect 14280 18702 14332 18708
rect 14464 18760 14516 18766
rect 14464 18702 14516 18708
rect 13740 17190 13860 17218
rect 13648 17088 13768 17116
rect 13360 17070 13412 17076
rect 12912 16658 12940 17070
rect 13268 17060 13320 17066
rect 13268 17002 13320 17008
rect 12900 16652 12952 16658
rect 12900 16594 12952 16600
rect 12992 16108 13044 16114
rect 12992 16050 13044 16056
rect 13004 15706 13032 16050
rect 13280 16046 13308 17002
rect 13636 16992 13688 16998
rect 13636 16934 13688 16940
rect 13360 16652 13412 16658
rect 13360 16594 13412 16600
rect 13084 16040 13136 16046
rect 13084 15982 13136 15988
rect 13268 16040 13320 16046
rect 13268 15982 13320 15988
rect 12992 15700 13044 15706
rect 12992 15642 13044 15648
rect 12452 13326 12480 13670
rect 12544 13654 12664 13682
rect 12440 13320 12492 13326
rect 12440 13262 12492 13268
rect 12256 12844 12308 12850
rect 12256 12786 12308 12792
rect 11244 12776 11296 12782
rect 11244 12718 11296 12724
rect 11152 12640 11204 12646
rect 11152 12582 11204 12588
rect 11060 12368 11112 12374
rect 11060 12310 11112 12316
rect 11164 12238 11192 12582
rect 11152 12232 11204 12238
rect 11152 12174 11204 12180
rect 10876 12096 10928 12102
rect 10876 12038 10928 12044
rect 10600 11688 10652 11694
rect 10600 11630 10652 11636
rect 10888 11082 10916 12038
rect 11256 11898 11284 12718
rect 12452 12306 12480 13262
rect 12636 13258 12664 13654
rect 12624 13252 12676 13258
rect 12624 13194 12676 13200
rect 12440 12300 12492 12306
rect 12440 12242 12492 12248
rect 11244 11892 11296 11898
rect 11244 11834 11296 11840
rect 11888 11892 11940 11898
rect 11888 11834 11940 11840
rect 11796 11688 11848 11694
rect 11796 11630 11848 11636
rect 11152 11552 11204 11558
rect 11152 11494 11204 11500
rect 10416 11076 10468 11082
rect 10416 11018 10468 11024
rect 10876 11076 10928 11082
rect 10876 11018 10928 11024
rect 10428 10810 10456 11018
rect 10140 10804 10192 10810
rect 10140 10746 10192 10752
rect 10232 10804 10284 10810
rect 10232 10746 10284 10752
rect 10416 10804 10468 10810
rect 10416 10746 10468 10752
rect 10244 9722 10272 10746
rect 11164 10674 11192 11494
rect 11808 10742 11836 11630
rect 11900 11354 11928 11834
rect 12636 11762 12664 13194
rect 12808 12912 12860 12918
rect 12808 12854 12860 12860
rect 12348 11756 12400 11762
rect 12348 11698 12400 11704
rect 12624 11756 12676 11762
rect 12624 11698 12676 11704
rect 12360 11354 12388 11698
rect 11888 11348 11940 11354
rect 11888 11290 11940 11296
rect 12348 11348 12400 11354
rect 12348 11290 12400 11296
rect 11796 10736 11848 10742
rect 11716 10696 11796 10724
rect 11152 10668 11204 10674
rect 11152 10610 11204 10616
rect 10784 9988 10836 9994
rect 10784 9930 10836 9936
rect 10232 9716 10284 9722
rect 10232 9658 10284 9664
rect 9772 9444 9824 9450
rect 9772 9386 9824 9392
rect 9864 9376 9916 9382
rect 9864 9318 9916 9324
rect 9876 8974 9904 9318
rect 10796 9178 10824 9930
rect 10876 9920 10928 9926
rect 10876 9862 10928 9868
rect 10888 9654 10916 9862
rect 10876 9648 10928 9654
rect 10876 9590 10928 9596
rect 11716 9586 11744 10696
rect 11796 10678 11848 10684
rect 11796 10600 11848 10606
rect 11796 10542 11848 10548
rect 11808 10266 11836 10542
rect 11796 10260 11848 10266
rect 11796 10202 11848 10208
rect 12072 9648 12124 9654
rect 12072 9590 12124 9596
rect 10968 9580 11020 9586
rect 10968 9522 11020 9528
rect 11704 9580 11756 9586
rect 11704 9522 11756 9528
rect 10980 9178 11008 9522
rect 10784 9172 10836 9178
rect 10784 9114 10836 9120
rect 10968 9172 11020 9178
rect 10968 9114 11020 9120
rect 9864 8968 9916 8974
rect 9864 8910 9916 8916
rect 10876 8832 10928 8838
rect 10876 8774 10928 8780
rect 10888 8566 10916 8774
rect 12084 8634 12112 9590
rect 12072 8628 12124 8634
rect 12072 8570 12124 8576
rect 10416 8560 10468 8566
rect 10416 8502 10468 8508
rect 10876 8560 10928 8566
rect 10876 8502 10928 8508
rect 12440 8560 12492 8566
rect 12440 8502 12492 8508
rect 9220 8424 9272 8430
rect 9220 8366 9272 8372
rect 8300 7948 8352 7954
rect 8300 7890 8352 7896
rect 8024 7812 8076 7818
rect 8024 7754 8076 7760
rect 8944 7744 8996 7750
rect 8944 7686 8996 7692
rect 9036 7744 9088 7750
rect 9036 7686 9088 7692
rect 8956 7478 8984 7686
rect 9048 7546 9076 7686
rect 9036 7540 9088 7546
rect 9036 7482 9088 7488
rect 8944 7472 8996 7478
rect 8944 7414 8996 7420
rect 9232 7410 9260 8366
rect 10428 8090 10456 8502
rect 11796 8424 11848 8430
rect 11796 8366 11848 8372
rect 10416 8084 10468 8090
rect 10416 8026 10468 8032
rect 11808 7410 11836 8366
rect 12452 7886 12480 8502
rect 12440 7880 12492 7886
rect 12440 7822 12492 7828
rect 12452 7410 12480 7822
rect 12636 7818 12664 11698
rect 12820 11218 12848 12854
rect 13096 12850 13124 15982
rect 13280 15570 13308 15982
rect 13268 15564 13320 15570
rect 13268 15506 13320 15512
rect 13372 15094 13400 16594
rect 13648 16590 13676 16934
rect 13740 16794 13768 17088
rect 13728 16788 13780 16794
rect 13728 16730 13780 16736
rect 13636 16584 13688 16590
rect 13636 16526 13688 16532
rect 13544 16448 13596 16454
rect 13544 16390 13596 16396
rect 13556 16182 13584 16390
rect 13832 16250 13860 17190
rect 14096 17196 14148 17202
rect 14096 17138 14148 17144
rect 14108 16726 14136 17138
rect 14096 16720 14148 16726
rect 14096 16662 14148 16668
rect 13820 16244 13872 16250
rect 13820 16186 13872 16192
rect 13544 16176 13596 16182
rect 13544 16118 13596 16124
rect 14108 16046 14136 16662
rect 14292 16658 14320 18702
rect 14476 18222 14504 18702
rect 14464 18216 14516 18222
rect 14464 18158 14516 18164
rect 14280 16652 14332 16658
rect 14280 16594 14332 16600
rect 14660 16590 14688 22646
rect 14844 22094 14872 28426
rect 14936 22710 14964 30194
rect 15568 30184 15620 30190
rect 15568 30126 15620 30132
rect 15292 30048 15344 30054
rect 15292 29990 15344 29996
rect 15304 29102 15332 29990
rect 15580 29850 15608 30126
rect 15764 29850 15792 30194
rect 16224 30190 16252 33390
rect 16684 32978 16712 33390
rect 16672 32972 16724 32978
rect 16672 32914 16724 32920
rect 16684 32366 16712 32914
rect 16868 32842 16896 33798
rect 16856 32836 16908 32842
rect 16856 32778 16908 32784
rect 16856 32428 16908 32434
rect 16856 32370 16908 32376
rect 16672 32360 16724 32366
rect 16672 32302 16724 32308
rect 16580 31136 16632 31142
rect 16580 31078 16632 31084
rect 16396 30660 16448 30666
rect 16396 30602 16448 30608
rect 16408 30326 16436 30602
rect 16592 30598 16620 31078
rect 16580 30592 16632 30598
rect 16580 30534 16632 30540
rect 16592 30394 16620 30534
rect 16580 30388 16632 30394
rect 16580 30330 16632 30336
rect 16396 30320 16448 30326
rect 16396 30262 16448 30268
rect 16212 30184 16264 30190
rect 16212 30126 16264 30132
rect 16868 30054 16896 32370
rect 17052 30258 17080 34070
rect 17144 33522 17172 36654
rect 17328 36106 17356 37062
rect 17972 36922 18000 37062
rect 17960 36916 18012 36922
rect 17960 36858 18012 36864
rect 18156 36378 18184 38150
rect 18616 38010 18644 38218
rect 18604 38004 18656 38010
rect 18604 37946 18656 37952
rect 18236 37868 18288 37874
rect 18236 37810 18288 37816
rect 18144 36372 18196 36378
rect 18144 36314 18196 36320
rect 18248 36310 18276 37810
rect 18708 37330 18736 38354
rect 19076 37874 19104 38422
rect 19260 38010 19288 38508
rect 22284 38490 22336 38496
rect 25228 38548 25280 38554
rect 25228 38490 25280 38496
rect 28184 38486 28212 40093
rect 30288 38548 30340 38554
rect 30288 38490 30340 38496
rect 28172 38480 28224 38486
rect 19984 38412 20036 38418
rect 19984 38354 20036 38360
rect 20352 38412 20404 38418
rect 20352 38354 20404 38360
rect 23492 38406 23704 38434
rect 28172 38422 28224 38428
rect 19524 38344 19576 38350
rect 19524 38286 19576 38292
rect 19432 38208 19484 38214
rect 19432 38150 19484 38156
rect 19248 38004 19300 38010
rect 19248 37946 19300 37952
rect 19064 37868 19116 37874
rect 19064 37810 19116 37816
rect 18696 37324 18748 37330
rect 18696 37266 18748 37272
rect 18328 37188 18380 37194
rect 18328 37130 18380 37136
rect 18340 36922 18368 37130
rect 18604 37120 18656 37126
rect 18604 37062 18656 37068
rect 18328 36916 18380 36922
rect 18328 36858 18380 36864
rect 18328 36780 18380 36786
rect 18328 36722 18380 36728
rect 18236 36304 18288 36310
rect 18236 36246 18288 36252
rect 18340 36174 18368 36722
rect 18616 36310 18644 37062
rect 18604 36304 18656 36310
rect 18604 36246 18656 36252
rect 17684 36168 17736 36174
rect 17684 36110 17736 36116
rect 17960 36168 18012 36174
rect 17960 36110 18012 36116
rect 18328 36168 18380 36174
rect 18328 36110 18380 36116
rect 17316 36100 17368 36106
rect 17316 36042 17368 36048
rect 17328 35154 17356 36042
rect 17696 35766 17724 36110
rect 17684 35760 17736 35766
rect 17684 35702 17736 35708
rect 17868 35692 17920 35698
rect 17868 35634 17920 35640
rect 17316 35148 17368 35154
rect 17316 35090 17368 35096
rect 17880 34746 17908 35634
rect 17972 35630 18000 36110
rect 17960 35624 18012 35630
rect 17960 35566 18012 35572
rect 17972 35290 18000 35566
rect 17960 35284 18012 35290
rect 17960 35226 18012 35232
rect 18616 34746 18644 36246
rect 18708 35630 18736 37266
rect 19444 37262 19472 38150
rect 19432 37256 19484 37262
rect 19432 37198 19484 37204
rect 19156 36848 19208 36854
rect 19156 36790 19208 36796
rect 19168 35834 19196 36790
rect 19432 36576 19484 36582
rect 19432 36518 19484 36524
rect 19444 36106 19472 36518
rect 19536 36174 19564 38286
rect 19892 38208 19944 38214
rect 19892 38150 19944 38156
rect 19904 37942 19932 38150
rect 19892 37936 19944 37942
rect 19892 37878 19944 37884
rect 19616 37664 19668 37670
rect 19616 37606 19668 37612
rect 19628 37262 19656 37606
rect 19616 37256 19668 37262
rect 19616 37198 19668 37204
rect 19708 37120 19760 37126
rect 19708 37062 19760 37068
rect 19720 36854 19748 37062
rect 19708 36848 19760 36854
rect 19708 36790 19760 36796
rect 19996 36242 20024 38354
rect 20364 37806 20392 38354
rect 23492 38350 23520 38406
rect 23676 38350 23704 38406
rect 29552 38412 29604 38418
rect 29552 38354 29604 38360
rect 22560 38344 22612 38350
rect 22560 38286 22612 38292
rect 23480 38344 23532 38350
rect 23480 38286 23532 38292
rect 23664 38344 23716 38350
rect 23664 38286 23716 38292
rect 24768 38344 24820 38350
rect 24768 38286 24820 38292
rect 25412 38344 25464 38350
rect 25412 38286 25464 38292
rect 28540 38344 28592 38350
rect 28540 38286 28592 38292
rect 21364 38208 21416 38214
rect 21364 38150 21416 38156
rect 21376 37874 21404 38150
rect 22008 37936 22060 37942
rect 22008 37878 22060 37884
rect 21364 37868 21416 37874
rect 21364 37810 21416 37816
rect 20168 37800 20220 37806
rect 20168 37742 20220 37748
rect 20352 37800 20404 37806
rect 20352 37742 20404 37748
rect 20180 37194 20208 37742
rect 20260 37256 20312 37262
rect 20260 37198 20312 37204
rect 20168 37188 20220 37194
rect 20168 37130 20220 37136
rect 19708 36236 19760 36242
rect 19708 36178 19760 36184
rect 19984 36236 20036 36242
rect 19984 36178 20036 36184
rect 19524 36168 19576 36174
rect 19524 36110 19576 36116
rect 19432 36100 19484 36106
rect 19432 36042 19484 36048
rect 19156 35828 19208 35834
rect 19156 35770 19208 35776
rect 19248 35692 19300 35698
rect 19248 35634 19300 35640
rect 18696 35624 18748 35630
rect 18696 35566 18748 35572
rect 19260 35086 19288 35634
rect 19248 35080 19300 35086
rect 19248 35022 19300 35028
rect 19340 34944 19392 34950
rect 19340 34886 19392 34892
rect 17868 34740 17920 34746
rect 17868 34682 17920 34688
rect 18604 34740 18656 34746
rect 18604 34682 18656 34688
rect 18052 34604 18104 34610
rect 18052 34546 18104 34552
rect 18420 34604 18472 34610
rect 18420 34546 18472 34552
rect 17868 34400 17920 34406
rect 17868 34342 17920 34348
rect 17408 33992 17460 33998
rect 17408 33934 17460 33940
rect 17132 33516 17184 33522
rect 17132 33458 17184 33464
rect 17420 33114 17448 33934
rect 17592 33856 17644 33862
rect 17592 33798 17644 33804
rect 17500 33652 17552 33658
rect 17500 33594 17552 33600
rect 17408 33108 17460 33114
rect 17408 33050 17460 33056
rect 17512 32774 17540 33594
rect 17604 33590 17632 33798
rect 17880 33590 17908 34342
rect 17592 33584 17644 33590
rect 17592 33526 17644 33532
rect 17868 33584 17920 33590
rect 17868 33526 17920 33532
rect 17960 32904 18012 32910
rect 17960 32846 18012 32852
rect 17500 32768 17552 32774
rect 17500 32710 17552 32716
rect 17868 32768 17920 32774
rect 17868 32710 17920 32716
rect 17132 32360 17184 32366
rect 17132 32302 17184 32308
rect 17144 31822 17172 32302
rect 17316 32224 17368 32230
rect 17316 32166 17368 32172
rect 17132 31816 17184 31822
rect 17132 31758 17184 31764
rect 17224 31408 17276 31414
rect 17224 31350 17276 31356
rect 17236 30326 17264 31350
rect 17328 30802 17356 32166
rect 17408 31748 17460 31754
rect 17408 31690 17460 31696
rect 17420 31482 17448 31690
rect 17684 31680 17736 31686
rect 17684 31622 17736 31628
rect 17776 31680 17828 31686
rect 17776 31622 17828 31628
rect 17408 31476 17460 31482
rect 17408 31418 17460 31424
rect 17316 30796 17368 30802
rect 17316 30738 17368 30744
rect 17696 30734 17724 31622
rect 17788 31414 17816 31622
rect 17776 31408 17828 31414
rect 17776 31350 17828 31356
rect 17880 31346 17908 32710
rect 17868 31340 17920 31346
rect 17868 31282 17920 31288
rect 17972 31142 18000 32846
rect 18064 32434 18092 34546
rect 18236 34400 18288 34406
rect 18236 34342 18288 34348
rect 18248 34202 18276 34342
rect 18236 34196 18288 34202
rect 18236 34138 18288 34144
rect 18432 33658 18460 34546
rect 19352 34066 19380 34886
rect 19444 34610 19472 36042
rect 19524 35624 19576 35630
rect 19524 35566 19576 35572
rect 19536 35018 19564 35566
rect 19524 35012 19576 35018
rect 19524 34954 19576 34960
rect 19432 34604 19484 34610
rect 19432 34546 19484 34552
rect 19340 34060 19392 34066
rect 19340 34002 19392 34008
rect 19064 33924 19116 33930
rect 19064 33866 19116 33872
rect 18880 33856 18932 33862
rect 18880 33798 18932 33804
rect 18420 33652 18472 33658
rect 18420 33594 18472 33600
rect 18432 32978 18460 33594
rect 18420 32972 18472 32978
rect 18420 32914 18472 32920
rect 18892 32842 18920 33798
rect 19076 33658 19104 33866
rect 19064 33652 19116 33658
rect 19064 33594 19116 33600
rect 19444 33590 19472 34546
rect 19432 33584 19484 33590
rect 19432 33526 19484 33532
rect 19536 33114 19564 34954
rect 19524 33108 19576 33114
rect 19524 33050 19576 33056
rect 18880 32836 18932 32842
rect 18880 32778 18932 32784
rect 18512 32768 18564 32774
rect 18512 32710 18564 32716
rect 18524 32570 18552 32710
rect 18512 32564 18564 32570
rect 18512 32506 18564 32512
rect 18052 32428 18104 32434
rect 18052 32370 18104 32376
rect 19524 32428 19576 32434
rect 19524 32370 19576 32376
rect 17960 31136 18012 31142
rect 17960 31078 18012 31084
rect 17684 30728 17736 30734
rect 17684 30670 17736 30676
rect 17696 30326 17724 30670
rect 17224 30320 17276 30326
rect 17224 30262 17276 30268
rect 17684 30320 17736 30326
rect 17684 30262 17736 30268
rect 18064 30258 18092 32370
rect 18512 32224 18564 32230
rect 18512 32166 18564 32172
rect 18524 31822 18552 32166
rect 19536 31890 19564 32370
rect 19720 32366 19748 36178
rect 20180 36174 20208 37130
rect 20272 36718 20300 37198
rect 20260 36712 20312 36718
rect 20260 36654 20312 36660
rect 20168 36168 20220 36174
rect 20168 36110 20220 36116
rect 19984 36032 20036 36038
rect 19984 35974 20036 35980
rect 19996 35894 20024 35974
rect 19812 35866 20024 35894
rect 19812 34950 19840 35866
rect 19892 35760 19944 35766
rect 19892 35702 19944 35708
rect 19904 35154 19932 35702
rect 20364 35154 20392 37742
rect 21272 37188 21324 37194
rect 21272 37130 21324 37136
rect 21284 36922 21312 37130
rect 22020 37126 22048 37878
rect 22572 37466 22600 38286
rect 23572 38276 23624 38282
rect 23572 38218 23624 38224
rect 23112 38208 23164 38214
rect 23112 38150 23164 38156
rect 22744 37936 22796 37942
rect 22744 37878 22796 37884
rect 22560 37460 22612 37466
rect 22560 37402 22612 37408
rect 22008 37120 22060 37126
rect 22006 37088 22008 37097
rect 22376 37120 22428 37126
rect 22060 37088 22062 37097
rect 22376 37062 22428 37068
rect 22006 37023 22062 37032
rect 22020 36997 22048 37023
rect 21272 36916 21324 36922
rect 21272 36858 21324 36864
rect 22388 36854 22416 37062
rect 22376 36848 22428 36854
rect 22376 36790 22428 36796
rect 21272 36780 21324 36786
rect 21272 36722 21324 36728
rect 21284 36106 21312 36722
rect 22100 36712 22152 36718
rect 22100 36654 22152 36660
rect 21272 36100 21324 36106
rect 21272 36042 21324 36048
rect 20444 36032 20496 36038
rect 20444 35974 20496 35980
rect 20456 35834 20484 35974
rect 20444 35828 20496 35834
rect 20444 35770 20496 35776
rect 20904 35488 20956 35494
rect 20904 35430 20956 35436
rect 19892 35148 19944 35154
rect 19892 35090 19944 35096
rect 19984 35148 20036 35154
rect 19984 35090 20036 35096
rect 20352 35148 20404 35154
rect 20352 35090 20404 35096
rect 19800 34944 19852 34950
rect 19800 34886 19852 34892
rect 19812 34542 19840 34886
rect 19800 34536 19852 34542
rect 19800 34478 19852 34484
rect 19996 34066 20024 35090
rect 20916 35018 20944 35430
rect 20904 35012 20956 35018
rect 20904 34954 20956 34960
rect 20812 34604 20864 34610
rect 20812 34546 20864 34552
rect 20824 34202 20852 34546
rect 20812 34196 20864 34202
rect 20812 34138 20864 34144
rect 19984 34060 20036 34066
rect 19984 34002 20036 34008
rect 19800 33856 19852 33862
rect 19800 33798 19852 33804
rect 19812 33114 19840 33798
rect 19800 33108 19852 33114
rect 19800 33050 19852 33056
rect 19812 32570 19840 33050
rect 19800 32564 19852 32570
rect 19800 32506 19852 32512
rect 19708 32360 19760 32366
rect 19708 32302 19760 32308
rect 19524 31884 19576 31890
rect 19524 31826 19576 31832
rect 18512 31816 18564 31822
rect 18512 31758 18564 31764
rect 19616 31816 19668 31822
rect 19616 31758 19668 31764
rect 19432 31680 19484 31686
rect 19432 31622 19484 31628
rect 19064 31476 19116 31482
rect 19064 31418 19116 31424
rect 18512 30728 18564 30734
rect 18512 30670 18564 30676
rect 18524 30258 18552 30670
rect 19076 30394 19104 31418
rect 19156 31272 19208 31278
rect 19156 31214 19208 31220
rect 19340 31272 19392 31278
rect 19340 31214 19392 31220
rect 19168 30734 19196 31214
rect 19352 30938 19380 31214
rect 19340 30932 19392 30938
rect 19340 30874 19392 30880
rect 19156 30728 19208 30734
rect 19156 30670 19208 30676
rect 19064 30388 19116 30394
rect 19064 30330 19116 30336
rect 19444 30326 19472 31622
rect 19628 30938 19656 31758
rect 19616 30932 19668 30938
rect 19616 30874 19668 30880
rect 19432 30320 19484 30326
rect 19432 30262 19484 30268
rect 17040 30252 17092 30258
rect 17040 30194 17092 30200
rect 18052 30252 18104 30258
rect 18052 30194 18104 30200
rect 18512 30252 18564 30258
rect 18512 30194 18564 30200
rect 16856 30048 16908 30054
rect 16856 29990 16908 29996
rect 15568 29844 15620 29850
rect 15568 29786 15620 29792
rect 15752 29844 15804 29850
rect 15752 29786 15804 29792
rect 18144 29708 18196 29714
rect 18144 29650 18196 29656
rect 17500 29640 17552 29646
rect 17500 29582 17552 29588
rect 15476 29572 15528 29578
rect 15476 29514 15528 29520
rect 15292 29096 15344 29102
rect 15292 29038 15344 29044
rect 15488 28558 15516 29514
rect 16120 29504 16172 29510
rect 16120 29446 16172 29452
rect 16304 29504 16356 29510
rect 16304 29446 16356 29452
rect 15568 29232 15620 29238
rect 15568 29174 15620 29180
rect 15580 28762 15608 29174
rect 16132 28762 16160 29446
rect 16316 28966 16344 29446
rect 16304 28960 16356 28966
rect 16304 28902 16356 28908
rect 15568 28756 15620 28762
rect 15568 28698 15620 28704
rect 16120 28756 16172 28762
rect 16120 28698 16172 28704
rect 15476 28552 15528 28558
rect 15476 28494 15528 28500
rect 16120 28416 16172 28422
rect 16120 28358 16172 28364
rect 15016 27940 15068 27946
rect 15016 27882 15068 27888
rect 15028 26926 15056 27882
rect 16132 27674 16160 28358
rect 16316 28150 16344 28902
rect 16856 28552 16908 28558
rect 16856 28494 16908 28500
rect 16868 28218 16896 28494
rect 16856 28212 16908 28218
rect 16856 28154 16908 28160
rect 16304 28144 16356 28150
rect 16304 28086 16356 28092
rect 16120 27668 16172 27674
rect 16120 27610 16172 27616
rect 16488 27328 16540 27334
rect 16488 27270 16540 27276
rect 15016 26920 15068 26926
rect 15016 26862 15068 26868
rect 15108 26852 15160 26858
rect 15108 26794 15160 26800
rect 15120 26450 15148 26794
rect 15108 26444 15160 26450
rect 15108 26386 15160 26392
rect 15200 25968 15252 25974
rect 15200 25910 15252 25916
rect 15212 24750 15240 25910
rect 15660 25832 15712 25838
rect 15660 25774 15712 25780
rect 15292 25220 15344 25226
rect 15292 25162 15344 25168
rect 15304 24818 15332 25162
rect 15292 24812 15344 24818
rect 15292 24754 15344 24760
rect 15200 24744 15252 24750
rect 15200 24686 15252 24692
rect 15672 24410 15700 25774
rect 16304 25696 16356 25702
rect 16304 25638 16356 25644
rect 16316 25362 16344 25638
rect 16304 25356 16356 25362
rect 16304 25298 16356 25304
rect 15936 25152 15988 25158
rect 15936 25094 15988 25100
rect 15660 24404 15712 24410
rect 15660 24346 15712 24352
rect 15476 24064 15528 24070
rect 15476 24006 15528 24012
rect 15200 23724 15252 23730
rect 15200 23666 15252 23672
rect 14924 22704 14976 22710
rect 14924 22646 14976 22652
rect 14924 22094 14976 22098
rect 14844 22092 14976 22094
rect 14844 22066 14924 22092
rect 14924 22034 14976 22040
rect 15016 21956 15068 21962
rect 15016 21898 15068 21904
rect 15028 21690 15056 21898
rect 15016 21684 15068 21690
rect 15016 21626 15068 21632
rect 14740 21412 14792 21418
rect 14740 21354 14792 21360
rect 14752 19990 14780 21354
rect 14740 19984 14792 19990
rect 14740 19926 14792 19932
rect 15212 18714 15240 23666
rect 15488 23186 15516 24006
rect 15476 23180 15528 23186
rect 15476 23122 15528 23128
rect 15568 22500 15620 22506
rect 15568 22442 15620 22448
rect 15580 22166 15608 22442
rect 15568 22160 15620 22166
rect 15568 22102 15620 22108
rect 15844 21548 15896 21554
rect 15844 21490 15896 21496
rect 15856 21146 15884 21490
rect 15844 21140 15896 21146
rect 15844 21082 15896 21088
rect 15384 20800 15436 20806
rect 15384 20742 15436 20748
rect 15660 20800 15712 20806
rect 15660 20742 15712 20748
rect 15396 20534 15424 20742
rect 15672 20602 15700 20742
rect 15660 20596 15712 20602
rect 15660 20538 15712 20544
rect 15384 20528 15436 20534
rect 15384 20470 15436 20476
rect 15660 19848 15712 19854
rect 15660 19790 15712 19796
rect 15672 19514 15700 19790
rect 15660 19508 15712 19514
rect 15660 19450 15712 19456
rect 15292 19440 15344 19446
rect 15292 19382 15344 19388
rect 15304 18970 15332 19382
rect 15292 18964 15344 18970
rect 15292 18906 15344 18912
rect 15660 18964 15712 18970
rect 15660 18906 15712 18912
rect 15212 18686 15332 18714
rect 14924 18624 14976 18630
rect 14924 18566 14976 18572
rect 15200 18624 15252 18630
rect 15200 18566 15252 18572
rect 14936 17678 14964 18566
rect 15212 18426 15240 18566
rect 15200 18420 15252 18426
rect 15200 18362 15252 18368
rect 15304 18306 15332 18686
rect 15476 18692 15528 18698
rect 15476 18634 15528 18640
rect 15212 18278 15332 18306
rect 14924 17672 14976 17678
rect 14924 17614 14976 17620
rect 14832 17128 14884 17134
rect 14832 17070 14884 17076
rect 14648 16584 14700 16590
rect 14648 16526 14700 16532
rect 14464 16516 14516 16522
rect 14464 16458 14516 16464
rect 14096 16040 14148 16046
rect 14096 15982 14148 15988
rect 13820 15632 13872 15638
rect 13820 15574 13872 15580
rect 13832 15094 13860 15574
rect 14476 15094 14504 16458
rect 13360 15088 13412 15094
rect 13360 15030 13412 15036
rect 13820 15088 13872 15094
rect 13820 15030 13872 15036
rect 14464 15088 14516 15094
rect 14464 15030 14516 15036
rect 13832 14414 13860 15030
rect 13820 14408 13872 14414
rect 13820 14350 13872 14356
rect 13820 14272 13872 14278
rect 13820 14214 13872 14220
rect 13832 14074 13860 14214
rect 13820 14068 13872 14074
rect 13820 14010 13872 14016
rect 13728 14000 13780 14006
rect 13728 13942 13780 13948
rect 13636 13932 13688 13938
rect 13636 13874 13688 13880
rect 13360 13864 13412 13870
rect 13360 13806 13412 13812
rect 13372 13190 13400 13806
rect 13360 13184 13412 13190
rect 13360 13126 13412 13132
rect 13544 12912 13596 12918
rect 13544 12854 13596 12860
rect 13084 12844 13136 12850
rect 13084 12786 13136 12792
rect 13556 12442 13584 12854
rect 13544 12436 13596 12442
rect 13544 12378 13596 12384
rect 13648 11830 13676 13874
rect 13740 12986 13768 13942
rect 14660 13326 14688 16526
rect 14844 15706 14872 17070
rect 15108 16176 15160 16182
rect 15108 16118 15160 16124
rect 14832 15700 14884 15706
rect 14832 15642 14884 15648
rect 15120 15162 15148 16118
rect 15212 15978 15240 18278
rect 15488 18222 15516 18634
rect 15292 18216 15344 18222
rect 15292 18158 15344 18164
rect 15476 18216 15528 18222
rect 15476 18158 15528 18164
rect 15304 17746 15332 18158
rect 15292 17740 15344 17746
rect 15292 17682 15344 17688
rect 15304 17134 15332 17682
rect 15384 17536 15436 17542
rect 15384 17478 15436 17484
rect 15292 17128 15344 17134
rect 15292 17070 15344 17076
rect 15200 15972 15252 15978
rect 15200 15914 15252 15920
rect 15212 15502 15240 15914
rect 15396 15502 15424 17478
rect 15568 17264 15620 17270
rect 15568 17206 15620 17212
rect 15580 16250 15608 17206
rect 15672 16590 15700 18906
rect 15660 16584 15712 16590
rect 15660 16526 15712 16532
rect 15568 16244 15620 16250
rect 15568 16186 15620 16192
rect 15200 15496 15252 15502
rect 15200 15438 15252 15444
rect 15384 15496 15436 15502
rect 15384 15438 15436 15444
rect 15384 15360 15436 15366
rect 15384 15302 15436 15308
rect 15108 15156 15160 15162
rect 15108 15098 15160 15104
rect 15396 15026 15424 15302
rect 14740 15020 14792 15026
rect 14740 14962 14792 14968
rect 15384 15020 15436 15026
rect 15384 14962 15436 14968
rect 13820 13320 13872 13326
rect 13820 13262 13872 13268
rect 14648 13320 14700 13326
rect 14648 13262 14700 13268
rect 13728 12980 13780 12986
rect 13728 12922 13780 12928
rect 13832 12850 13860 13262
rect 14188 13184 14240 13190
rect 14188 13126 14240 13132
rect 13820 12844 13872 12850
rect 13820 12786 13872 12792
rect 14200 12714 14228 13126
rect 14660 12850 14688 13262
rect 14464 12844 14516 12850
rect 14464 12786 14516 12792
rect 14648 12844 14700 12850
rect 14648 12786 14700 12792
rect 14188 12708 14240 12714
rect 14188 12650 14240 12656
rect 13636 11824 13688 11830
rect 13636 11766 13688 11772
rect 12808 11212 12860 11218
rect 12808 11154 12860 11160
rect 13544 11076 13596 11082
rect 13544 11018 13596 11024
rect 12716 11008 12768 11014
rect 12716 10950 12768 10956
rect 12728 10130 12756 10950
rect 13556 10674 13584 11018
rect 13544 10668 13596 10674
rect 13544 10610 13596 10616
rect 12716 10124 12768 10130
rect 13648 10112 13676 11766
rect 13912 10464 13964 10470
rect 13912 10406 13964 10412
rect 12716 10066 12768 10072
rect 13556 10084 13676 10112
rect 12728 9722 12756 10066
rect 12716 9716 12768 9722
rect 12716 9658 12768 9664
rect 12728 8906 12756 9658
rect 13556 8974 13584 10084
rect 13924 10062 13952 10406
rect 13912 10056 13964 10062
rect 13912 9998 13964 10004
rect 13924 9722 13952 9998
rect 13912 9716 13964 9722
rect 13912 9658 13964 9664
rect 13912 9376 13964 9382
rect 13912 9318 13964 9324
rect 13924 9042 13952 9318
rect 14200 9110 14228 12650
rect 14476 12238 14504 12786
rect 14464 12232 14516 12238
rect 14464 12174 14516 12180
rect 14476 11150 14504 12174
rect 14752 11762 14780 14962
rect 15856 14958 15884 21082
rect 15948 20602 15976 25094
rect 16212 23520 16264 23526
rect 16212 23462 16264 23468
rect 16028 21888 16080 21894
rect 16028 21830 16080 21836
rect 16040 21622 16068 21830
rect 16028 21616 16080 21622
rect 16028 21558 16080 21564
rect 15936 20596 15988 20602
rect 15936 20538 15988 20544
rect 15948 19922 15976 20538
rect 16028 19984 16080 19990
rect 16028 19926 16080 19932
rect 15936 19916 15988 19922
rect 15936 19858 15988 19864
rect 16040 17814 16068 19926
rect 16224 18834 16252 23462
rect 16500 21486 16528 27270
rect 16764 27056 16816 27062
rect 16764 26998 16816 27004
rect 16580 25696 16632 25702
rect 16580 25638 16632 25644
rect 16592 23866 16620 25638
rect 16776 24750 16804 26998
rect 17408 26852 17460 26858
rect 17408 26794 17460 26800
rect 17224 26784 17276 26790
rect 17224 26726 17276 26732
rect 17236 25906 17264 26726
rect 17420 26450 17448 26794
rect 17408 26444 17460 26450
rect 17408 26386 17460 26392
rect 17224 25900 17276 25906
rect 17224 25842 17276 25848
rect 16948 25220 17000 25226
rect 16948 25162 17000 25168
rect 16764 24744 16816 24750
rect 16764 24686 16816 24692
rect 16672 24132 16724 24138
rect 16672 24074 16724 24080
rect 16684 23866 16712 24074
rect 16580 23860 16632 23866
rect 16580 23802 16632 23808
rect 16672 23860 16724 23866
rect 16672 23802 16724 23808
rect 16776 23730 16804 24686
rect 16960 24410 16988 25162
rect 17132 24608 17184 24614
rect 17132 24550 17184 24556
rect 16948 24404 17000 24410
rect 16948 24346 17000 24352
rect 17144 24274 17172 24550
rect 17132 24268 17184 24274
rect 17132 24210 17184 24216
rect 16764 23724 16816 23730
rect 16764 23666 16816 23672
rect 16776 23118 16804 23666
rect 17512 23118 17540 29582
rect 18156 28694 18184 29650
rect 18524 29646 18552 30194
rect 19720 29850 19748 32302
rect 19892 31884 19944 31890
rect 19892 31826 19944 31832
rect 19904 31346 19932 31826
rect 19892 31340 19944 31346
rect 19892 31282 19944 31288
rect 19904 30802 19932 31282
rect 19996 30802 20024 34002
rect 21284 33998 21312 36042
rect 21364 35692 21416 35698
rect 21364 35634 21416 35640
rect 21376 35290 21404 35634
rect 22008 35488 22060 35494
rect 22008 35430 22060 35436
rect 21364 35284 21416 35290
rect 21364 35226 21416 35232
rect 21376 33998 21404 35226
rect 22020 35086 22048 35430
rect 22112 35154 22140 36654
rect 22756 36378 22784 37878
rect 23020 37256 23072 37262
rect 23020 37198 23072 37204
rect 23032 36378 23060 37198
rect 23124 36854 23152 38150
rect 23584 37806 23612 38218
rect 23676 37890 23704 38286
rect 23756 38208 23808 38214
rect 23756 38150 23808 38156
rect 24492 38208 24544 38214
rect 24492 38150 24544 38156
rect 23768 38010 23796 38150
rect 23756 38004 23808 38010
rect 23756 37946 23808 37952
rect 24504 37942 24532 38150
rect 24492 37936 24544 37942
rect 23676 37862 23796 37890
rect 24492 37878 24544 37884
rect 23572 37800 23624 37806
rect 23572 37742 23624 37748
rect 23572 37324 23624 37330
rect 23572 37266 23624 37272
rect 23112 36848 23164 36854
rect 23112 36790 23164 36796
rect 23480 36576 23532 36582
rect 23480 36518 23532 36524
rect 22744 36372 22796 36378
rect 22744 36314 22796 36320
rect 23020 36372 23072 36378
rect 23020 36314 23072 36320
rect 23492 36242 23520 36518
rect 23584 36242 23612 37266
rect 23664 37120 23716 37126
rect 23664 37062 23716 37068
rect 23676 36922 23704 37062
rect 23664 36916 23716 36922
rect 23664 36858 23716 36864
rect 23480 36236 23532 36242
rect 23480 36178 23532 36184
rect 23572 36236 23624 36242
rect 23572 36178 23624 36184
rect 23388 36032 23440 36038
rect 23388 35974 23440 35980
rect 23400 35834 23428 35974
rect 23388 35828 23440 35834
rect 23388 35770 23440 35776
rect 22376 35760 22428 35766
rect 22376 35702 22428 35708
rect 22388 35290 22416 35702
rect 23296 35692 23348 35698
rect 23296 35634 23348 35640
rect 22744 35488 22796 35494
rect 22744 35430 22796 35436
rect 22376 35284 22428 35290
rect 22376 35226 22428 35232
rect 22192 35216 22244 35222
rect 22192 35158 22244 35164
rect 22100 35148 22152 35154
rect 22100 35090 22152 35096
rect 22008 35080 22060 35086
rect 22008 35022 22060 35028
rect 22112 34542 22140 35090
rect 22100 34536 22152 34542
rect 22100 34478 22152 34484
rect 20904 33992 20956 33998
rect 20904 33934 20956 33940
rect 21272 33992 21324 33998
rect 21272 33934 21324 33940
rect 21364 33992 21416 33998
rect 21364 33934 21416 33940
rect 20720 33516 20772 33522
rect 20720 33458 20772 33464
rect 20444 32836 20496 32842
rect 20444 32778 20496 32784
rect 20456 32570 20484 32778
rect 20444 32564 20496 32570
rect 20444 32506 20496 32512
rect 20076 32360 20128 32366
rect 20076 32302 20128 32308
rect 20088 31822 20116 32302
rect 20076 31816 20128 31822
rect 20076 31758 20128 31764
rect 20352 31816 20404 31822
rect 20352 31758 20404 31764
rect 19892 30796 19944 30802
rect 19892 30738 19944 30744
rect 19984 30796 20036 30802
rect 19984 30738 20036 30744
rect 19996 30190 20024 30738
rect 20364 30326 20392 31758
rect 20352 30320 20404 30326
rect 20352 30262 20404 30268
rect 19984 30184 20036 30190
rect 19984 30126 20036 30132
rect 19708 29844 19760 29850
rect 19708 29786 19760 29792
rect 18512 29640 18564 29646
rect 18512 29582 18564 29588
rect 18604 29640 18656 29646
rect 18604 29582 18656 29588
rect 18420 29504 18472 29510
rect 18420 29446 18472 29452
rect 18512 29504 18564 29510
rect 18512 29446 18564 29452
rect 18432 29306 18460 29446
rect 18420 29300 18472 29306
rect 18420 29242 18472 29248
rect 18144 28688 18196 28694
rect 18144 28630 18196 28636
rect 17592 28416 17644 28422
rect 17592 28358 17644 28364
rect 18052 28416 18104 28422
rect 18052 28358 18104 28364
rect 17604 28082 17632 28358
rect 18064 28082 18092 28358
rect 17592 28076 17644 28082
rect 17592 28018 17644 28024
rect 18052 28076 18104 28082
rect 18052 28018 18104 28024
rect 17604 27334 17632 28018
rect 17592 27328 17644 27334
rect 17592 27270 17644 27276
rect 17604 26382 17632 27270
rect 18156 26432 18184 28630
rect 18432 28626 18460 29242
rect 18236 28620 18288 28626
rect 18236 28562 18288 28568
rect 18420 28620 18472 28626
rect 18420 28562 18472 28568
rect 18248 27946 18276 28562
rect 18420 28416 18472 28422
rect 18420 28358 18472 28364
rect 18236 27940 18288 27946
rect 18236 27882 18288 27888
rect 18248 27538 18276 27882
rect 18432 27538 18460 28358
rect 18524 27606 18552 29446
rect 18616 29102 18644 29582
rect 19616 29572 19668 29578
rect 19616 29514 19668 29520
rect 19628 29170 19656 29514
rect 20260 29504 20312 29510
rect 20260 29446 20312 29452
rect 20272 29170 20300 29446
rect 19616 29164 19668 29170
rect 19616 29106 19668 29112
rect 20260 29164 20312 29170
rect 20260 29106 20312 29112
rect 18604 29096 18656 29102
rect 18604 29038 18656 29044
rect 18972 29096 19024 29102
rect 18972 29038 19024 29044
rect 18984 28626 19012 29038
rect 18696 28620 18748 28626
rect 18696 28562 18748 28568
rect 18972 28620 19024 28626
rect 18972 28562 19024 28568
rect 18708 28150 18736 28562
rect 18696 28144 18748 28150
rect 18696 28086 18748 28092
rect 18984 27878 19012 28562
rect 19892 28552 19944 28558
rect 19892 28494 19944 28500
rect 18972 27872 19024 27878
rect 18972 27814 19024 27820
rect 19708 27872 19760 27878
rect 19708 27814 19760 27820
rect 18512 27600 18564 27606
rect 18512 27542 18564 27548
rect 18236 27532 18288 27538
rect 18236 27474 18288 27480
rect 18420 27532 18472 27538
rect 18420 27474 18472 27480
rect 19340 27464 19392 27470
rect 19340 27406 19392 27412
rect 18880 27396 18932 27402
rect 18880 27338 18932 27344
rect 18420 27328 18472 27334
rect 18420 27270 18472 27276
rect 18432 26790 18460 27270
rect 18420 26784 18472 26790
rect 18420 26726 18472 26732
rect 18328 26580 18380 26586
rect 18328 26522 18380 26528
rect 18236 26444 18288 26450
rect 18156 26404 18236 26432
rect 18236 26386 18288 26392
rect 17592 26376 17644 26382
rect 17592 26318 17644 26324
rect 17960 25288 18012 25294
rect 17960 25230 18012 25236
rect 17868 24812 17920 24818
rect 17868 24754 17920 24760
rect 17880 24342 17908 24754
rect 17972 24682 18000 25230
rect 18248 24750 18276 26386
rect 18340 25974 18368 26522
rect 18432 26450 18460 26726
rect 18892 26586 18920 27338
rect 18972 26920 19024 26926
rect 18972 26862 19024 26868
rect 18984 26586 19012 26862
rect 18880 26580 18932 26586
rect 18880 26522 18932 26528
rect 18972 26580 19024 26586
rect 18972 26522 19024 26528
rect 18420 26444 18472 26450
rect 18420 26386 18472 26392
rect 18512 26240 18564 26246
rect 18512 26182 18564 26188
rect 18328 25968 18380 25974
rect 18328 25910 18380 25916
rect 18524 25498 18552 26182
rect 18604 25832 18656 25838
rect 18604 25774 18656 25780
rect 18512 25492 18564 25498
rect 18512 25434 18564 25440
rect 18052 24744 18104 24750
rect 18052 24686 18104 24692
rect 18236 24744 18288 24750
rect 18236 24686 18288 24692
rect 17960 24676 18012 24682
rect 17960 24618 18012 24624
rect 17868 24336 17920 24342
rect 17868 24278 17920 24284
rect 17776 24064 17828 24070
rect 17776 24006 17828 24012
rect 17788 23798 17816 24006
rect 17880 23866 17908 24278
rect 17868 23860 17920 23866
rect 17868 23802 17920 23808
rect 17776 23792 17828 23798
rect 17776 23734 17828 23740
rect 17592 23180 17644 23186
rect 17592 23122 17644 23128
rect 16764 23112 16816 23118
rect 16764 23054 16816 23060
rect 17500 23112 17552 23118
rect 17500 23054 17552 23060
rect 17316 22976 17368 22982
rect 17316 22918 17368 22924
rect 17328 22710 17356 22918
rect 17316 22704 17368 22710
rect 17316 22646 17368 22652
rect 17512 22030 17540 23054
rect 17604 22438 17632 23122
rect 17960 23112 18012 23118
rect 17960 23054 18012 23060
rect 17592 22432 17644 22438
rect 17592 22374 17644 22380
rect 17500 22024 17552 22030
rect 17500 21966 17552 21972
rect 17132 21956 17184 21962
rect 17132 21898 17184 21904
rect 16672 21888 16724 21894
rect 16672 21830 16724 21836
rect 16488 21480 16540 21486
rect 16488 21422 16540 21428
rect 16500 21350 16528 21422
rect 16488 21344 16540 21350
rect 16488 21286 16540 21292
rect 16684 20874 16712 21830
rect 16672 20868 16724 20874
rect 16672 20810 16724 20816
rect 16488 19236 16540 19242
rect 16488 19178 16540 19184
rect 16212 18828 16264 18834
rect 16212 18770 16264 18776
rect 16500 18766 16528 19178
rect 16580 18896 16632 18902
rect 16580 18838 16632 18844
rect 16488 18760 16540 18766
rect 16488 18702 16540 18708
rect 16592 18630 16620 18838
rect 16948 18828 17000 18834
rect 16948 18770 17000 18776
rect 16580 18624 16632 18630
rect 16580 18566 16632 18572
rect 16580 18352 16632 18358
rect 16580 18294 16632 18300
rect 16028 17808 16080 17814
rect 16028 17750 16080 17756
rect 16304 17604 16356 17610
rect 16304 17546 16356 17552
rect 16316 15094 16344 17546
rect 16488 17536 16540 17542
rect 16488 17478 16540 17484
rect 16500 17134 16528 17478
rect 16488 17128 16540 17134
rect 16488 17070 16540 17076
rect 16592 16522 16620 18294
rect 16764 18216 16816 18222
rect 16764 18158 16816 18164
rect 16776 17066 16804 18158
rect 16960 17746 16988 18770
rect 16948 17740 17000 17746
rect 16948 17682 17000 17688
rect 17144 17610 17172 21898
rect 17512 21622 17540 21966
rect 17500 21616 17552 21622
rect 17500 21558 17552 21564
rect 17604 21026 17632 22374
rect 17684 22228 17736 22234
rect 17684 22170 17736 22176
rect 17696 22098 17724 22170
rect 17684 22092 17736 22098
rect 17684 22034 17736 22040
rect 17776 21548 17828 21554
rect 17776 21490 17828 21496
rect 17604 20998 17724 21026
rect 17696 20942 17724 20998
rect 17684 20936 17736 20942
rect 17684 20878 17736 20884
rect 17408 20868 17460 20874
rect 17408 20810 17460 20816
rect 17420 20602 17448 20810
rect 17408 20596 17460 20602
rect 17408 20538 17460 20544
rect 17592 20256 17644 20262
rect 17592 20198 17644 20204
rect 17604 19786 17632 20198
rect 17696 19990 17724 20878
rect 17788 20806 17816 21490
rect 17972 21486 18000 23054
rect 17960 21480 18012 21486
rect 17960 21422 18012 21428
rect 18064 20874 18092 24686
rect 18328 24608 18380 24614
rect 18328 24550 18380 24556
rect 18340 24206 18368 24550
rect 18616 24206 18644 25774
rect 19352 25430 19380 27406
rect 19432 27328 19484 27334
rect 19432 27270 19484 27276
rect 19444 25770 19472 27270
rect 19720 26926 19748 27814
rect 19708 26920 19760 26926
rect 19708 26862 19760 26868
rect 19616 26784 19668 26790
rect 19616 26726 19668 26732
rect 19524 26240 19576 26246
rect 19524 26182 19576 26188
rect 19536 25906 19564 26182
rect 19524 25900 19576 25906
rect 19524 25842 19576 25848
rect 19432 25764 19484 25770
rect 19432 25706 19484 25712
rect 19340 25424 19392 25430
rect 19340 25366 19392 25372
rect 19064 24880 19116 24886
rect 19064 24822 19116 24828
rect 18972 24744 19024 24750
rect 18972 24686 19024 24692
rect 18328 24200 18380 24206
rect 18328 24142 18380 24148
rect 18604 24200 18656 24206
rect 18604 24142 18656 24148
rect 18512 23792 18564 23798
rect 18512 23734 18564 23740
rect 18524 23322 18552 23734
rect 18512 23316 18564 23322
rect 18512 23258 18564 23264
rect 18616 22642 18644 24142
rect 18604 22636 18656 22642
rect 18604 22578 18656 22584
rect 18616 22438 18644 22578
rect 18604 22432 18656 22438
rect 18604 22374 18656 22380
rect 18984 22166 19012 24686
rect 19076 23322 19104 24822
rect 19628 24274 19656 26726
rect 19720 26042 19748 26862
rect 19800 26852 19852 26858
rect 19800 26794 19852 26800
rect 19812 26518 19840 26794
rect 19904 26790 19932 28494
rect 19984 28416 20036 28422
rect 19984 28358 20036 28364
rect 20536 28416 20588 28422
rect 20536 28358 20588 28364
rect 19996 28150 20024 28358
rect 19984 28144 20036 28150
rect 19984 28086 20036 28092
rect 20444 27872 20496 27878
rect 20444 27814 20496 27820
rect 20456 27606 20484 27814
rect 20444 27600 20496 27606
rect 20444 27542 20496 27548
rect 20076 26988 20128 26994
rect 20076 26930 20128 26936
rect 19892 26784 19944 26790
rect 19892 26726 19944 26732
rect 19904 26518 19932 26726
rect 19800 26512 19852 26518
rect 19800 26454 19852 26460
rect 19892 26512 19944 26518
rect 19892 26454 19944 26460
rect 19892 26240 19944 26246
rect 19892 26182 19944 26188
rect 19708 26036 19760 26042
rect 19708 25978 19760 25984
rect 19720 25838 19748 25978
rect 19708 25832 19760 25838
rect 19708 25774 19760 25780
rect 19616 24268 19668 24274
rect 19616 24210 19668 24216
rect 19628 23322 19656 24210
rect 19720 23662 19748 25774
rect 19904 25684 19932 26182
rect 19984 25696 20036 25702
rect 19904 25656 19984 25684
rect 19904 25362 19932 25656
rect 19984 25638 20036 25644
rect 19892 25356 19944 25362
rect 19892 25298 19944 25304
rect 19800 25152 19852 25158
rect 19800 25094 19852 25100
rect 19812 24818 19840 25094
rect 19800 24812 19852 24818
rect 19800 24754 19852 24760
rect 19812 24274 19840 24754
rect 19984 24608 20036 24614
rect 19984 24550 20036 24556
rect 19800 24268 19852 24274
rect 19800 24210 19852 24216
rect 19812 23866 19840 24210
rect 19892 24064 19944 24070
rect 19892 24006 19944 24012
rect 19800 23860 19852 23866
rect 19800 23802 19852 23808
rect 19708 23656 19760 23662
rect 19708 23598 19760 23604
rect 19064 23316 19116 23322
rect 19064 23258 19116 23264
rect 19616 23316 19668 23322
rect 19616 23258 19668 23264
rect 19248 23112 19300 23118
rect 19248 23054 19300 23060
rect 19260 22642 19288 23054
rect 19248 22636 19300 22642
rect 19248 22578 19300 22584
rect 19248 22432 19300 22438
rect 19248 22374 19300 22380
rect 18972 22160 19024 22166
rect 18972 22102 19024 22108
rect 18236 22024 18288 22030
rect 18236 21966 18288 21972
rect 18248 21690 18276 21966
rect 18696 21888 18748 21894
rect 18696 21830 18748 21836
rect 18880 21888 18932 21894
rect 18880 21830 18932 21836
rect 18708 21690 18736 21830
rect 18236 21684 18288 21690
rect 18236 21626 18288 21632
rect 18696 21684 18748 21690
rect 18696 21626 18748 21632
rect 18236 21480 18288 21486
rect 18236 21422 18288 21428
rect 18052 20868 18104 20874
rect 18052 20810 18104 20816
rect 17776 20800 17828 20806
rect 17776 20742 17828 20748
rect 17788 20466 17816 20742
rect 17776 20460 17828 20466
rect 17776 20402 17828 20408
rect 17684 19984 17736 19990
rect 17684 19926 17736 19932
rect 17592 19780 17644 19786
rect 17592 19722 17644 19728
rect 17316 19304 17368 19310
rect 17316 19246 17368 19252
rect 17328 18766 17356 19246
rect 17788 18766 17816 20402
rect 17960 19712 18012 19718
rect 17960 19654 18012 19660
rect 17316 18760 17368 18766
rect 17316 18702 17368 18708
rect 17776 18760 17828 18766
rect 17776 18702 17828 18708
rect 17328 18086 17356 18702
rect 17500 18624 17552 18630
rect 17500 18566 17552 18572
rect 17316 18080 17368 18086
rect 17316 18022 17368 18028
rect 17328 17746 17356 18022
rect 17316 17740 17368 17746
rect 17316 17682 17368 17688
rect 17512 17610 17540 18566
rect 17132 17604 17184 17610
rect 17132 17546 17184 17552
rect 17500 17604 17552 17610
rect 17500 17546 17552 17552
rect 17512 17270 17540 17546
rect 17592 17536 17644 17542
rect 17592 17478 17644 17484
rect 17604 17338 17632 17478
rect 17592 17332 17644 17338
rect 17592 17274 17644 17280
rect 17500 17264 17552 17270
rect 17500 17206 17552 17212
rect 16764 17060 16816 17066
rect 16764 17002 16816 17008
rect 16776 16658 16804 17002
rect 16948 16992 17000 16998
rect 16948 16934 17000 16940
rect 16764 16652 16816 16658
rect 16764 16594 16816 16600
rect 16580 16516 16632 16522
rect 16580 16458 16632 16464
rect 16960 16114 16988 16934
rect 17132 16516 17184 16522
rect 17132 16458 17184 16464
rect 17144 16250 17172 16458
rect 17132 16244 17184 16250
rect 17132 16186 17184 16192
rect 16948 16108 17000 16114
rect 16948 16050 17000 16056
rect 17972 16046 18000 19654
rect 18052 19168 18104 19174
rect 18052 19110 18104 19116
rect 18064 17882 18092 19110
rect 18144 18352 18196 18358
rect 18144 18294 18196 18300
rect 18052 17876 18104 17882
rect 18052 17818 18104 17824
rect 18156 16810 18184 18294
rect 18064 16782 18184 16810
rect 18064 16454 18092 16782
rect 18144 16516 18196 16522
rect 18144 16458 18196 16464
rect 18052 16448 18104 16454
rect 18052 16390 18104 16396
rect 18156 16250 18184 16458
rect 18144 16244 18196 16250
rect 18144 16186 18196 16192
rect 18248 16182 18276 21422
rect 18696 21344 18748 21350
rect 18696 21286 18748 21292
rect 18512 20868 18564 20874
rect 18512 20810 18564 20816
rect 18236 16176 18288 16182
rect 18236 16118 18288 16124
rect 17960 16040 18012 16046
rect 17960 15982 18012 15988
rect 18524 15502 18552 20810
rect 18708 19854 18736 21286
rect 18892 19854 18920 21830
rect 19260 21622 19288 22374
rect 19720 22094 19748 23598
rect 19904 23186 19932 24006
rect 19996 23798 20024 24550
rect 19984 23792 20036 23798
rect 19984 23734 20036 23740
rect 19892 23180 19944 23186
rect 19892 23122 19944 23128
rect 19892 22976 19944 22982
rect 19892 22918 19944 22924
rect 19904 22574 19932 22918
rect 19892 22568 19944 22574
rect 19892 22510 19944 22516
rect 19904 22166 19932 22510
rect 19892 22160 19944 22166
rect 19892 22102 19944 22108
rect 19800 22094 19852 22098
rect 19720 22092 19852 22094
rect 19720 22066 19800 22092
rect 19800 22034 19852 22040
rect 19812 21622 19840 22034
rect 19248 21616 19300 21622
rect 19248 21558 19300 21564
rect 19800 21616 19852 21622
rect 19800 21558 19852 21564
rect 19708 21480 19760 21486
rect 19708 21422 19760 21428
rect 19432 20596 19484 20602
rect 19432 20538 19484 20544
rect 19156 20256 19208 20262
rect 19156 20198 19208 20204
rect 18696 19848 18748 19854
rect 18696 19790 18748 19796
rect 18880 19848 18932 19854
rect 18880 19790 18932 19796
rect 18788 19712 18840 19718
rect 18788 19654 18840 19660
rect 18972 19712 19024 19718
rect 18972 19654 19024 19660
rect 18800 18698 18828 19654
rect 18984 19514 19012 19654
rect 18972 19508 19024 19514
rect 18972 19450 19024 19456
rect 18880 19440 18932 19446
rect 18880 19382 18932 19388
rect 18892 18970 18920 19382
rect 19168 19310 19196 20198
rect 19156 19304 19208 19310
rect 19156 19246 19208 19252
rect 19444 18970 19472 20538
rect 19720 20058 19748 21422
rect 20088 21010 20116 26930
rect 20548 26330 20576 28358
rect 20628 27328 20680 27334
rect 20628 27270 20680 27276
rect 20640 27062 20668 27270
rect 20628 27056 20680 27062
rect 20628 26998 20680 27004
rect 20732 26994 20760 33458
rect 20916 32366 20944 33934
rect 21376 33810 21404 33934
rect 21284 33782 21404 33810
rect 21284 32434 21312 33782
rect 22112 33658 22140 34478
rect 22204 34406 22232 35158
rect 22756 34678 22784 35430
rect 23308 35290 23336 35634
rect 23296 35284 23348 35290
rect 23296 35226 23348 35232
rect 23584 35154 23612 36178
rect 23768 35630 23796 37862
rect 24216 37868 24268 37874
rect 24216 37810 24268 37816
rect 24228 37330 24256 37810
rect 24780 37466 24808 38286
rect 25228 38208 25280 38214
rect 25228 38150 25280 38156
rect 24768 37460 24820 37466
rect 24768 37402 24820 37408
rect 25240 37330 25268 38150
rect 24216 37324 24268 37330
rect 24216 37266 24268 37272
rect 24860 37324 24912 37330
rect 24860 37266 24912 37272
rect 25228 37324 25280 37330
rect 25228 37266 25280 37272
rect 24398 37088 24454 37097
rect 24398 37023 24454 37032
rect 24412 36922 24440 37023
rect 24400 36916 24452 36922
rect 24400 36858 24452 36864
rect 24032 36576 24084 36582
rect 24032 36518 24084 36524
rect 24044 35630 24072 36518
rect 24872 35698 24900 37266
rect 24952 36712 25004 36718
rect 24952 36654 25004 36660
rect 24964 36242 24992 36654
rect 25424 36650 25452 38286
rect 27712 38208 27764 38214
rect 27712 38150 27764 38156
rect 26424 37868 26476 37874
rect 26424 37810 26476 37816
rect 27160 37868 27212 37874
rect 27160 37810 27212 37816
rect 25504 37664 25556 37670
rect 25504 37606 25556 37612
rect 25516 37194 25544 37606
rect 25504 37188 25556 37194
rect 25504 37130 25556 37136
rect 25516 36786 25544 37130
rect 25504 36780 25556 36786
rect 25504 36722 25556 36728
rect 26148 36780 26200 36786
rect 26148 36722 26200 36728
rect 25412 36644 25464 36650
rect 25412 36586 25464 36592
rect 24952 36236 25004 36242
rect 24952 36178 25004 36184
rect 24964 36122 24992 36178
rect 24964 36094 25084 36122
rect 24952 36032 25004 36038
rect 24952 35974 25004 35980
rect 24964 35834 24992 35974
rect 24952 35828 25004 35834
rect 24952 35770 25004 35776
rect 24860 35692 24912 35698
rect 24860 35634 24912 35640
rect 23756 35624 23808 35630
rect 23756 35566 23808 35572
rect 24032 35624 24084 35630
rect 24032 35566 24084 35572
rect 23388 35148 23440 35154
rect 23388 35090 23440 35096
rect 23572 35148 23624 35154
rect 23572 35090 23624 35096
rect 23400 34950 23428 35090
rect 23388 34944 23440 34950
rect 23388 34886 23440 34892
rect 22744 34672 22796 34678
rect 22744 34614 22796 34620
rect 22192 34400 22244 34406
rect 22192 34342 22244 34348
rect 23400 34066 23428 34886
rect 23768 34610 23796 35566
rect 23940 34944 23992 34950
rect 23940 34886 23992 34892
rect 23952 34746 23980 34886
rect 23940 34740 23992 34746
rect 23940 34682 23992 34688
rect 24044 34626 24072 35566
rect 23756 34604 23808 34610
rect 23756 34546 23808 34552
rect 23952 34598 24072 34626
rect 23952 34542 23980 34598
rect 23940 34536 23992 34542
rect 23940 34478 23992 34484
rect 23388 34060 23440 34066
rect 23388 34002 23440 34008
rect 22284 33856 22336 33862
rect 22284 33798 22336 33804
rect 22836 33856 22888 33862
rect 22836 33798 22888 33804
rect 23848 33856 23900 33862
rect 23848 33798 23900 33804
rect 22100 33652 22152 33658
rect 22100 33594 22152 33600
rect 21824 33516 21876 33522
rect 21824 33458 21876 33464
rect 21836 32910 21864 33458
rect 22112 32978 22140 33594
rect 22296 33590 22324 33798
rect 22284 33584 22336 33590
rect 22284 33526 22336 33532
rect 22284 33448 22336 33454
rect 22284 33390 22336 33396
rect 22100 32972 22152 32978
rect 22100 32914 22152 32920
rect 21824 32904 21876 32910
rect 21824 32846 21876 32852
rect 21272 32428 21324 32434
rect 21272 32370 21324 32376
rect 20904 32360 20956 32366
rect 20904 32302 20956 32308
rect 21284 31346 21312 32370
rect 21456 32224 21508 32230
rect 21456 32166 21508 32172
rect 22008 32224 22060 32230
rect 22008 32166 22060 32172
rect 21468 31754 21496 32166
rect 22020 32026 22048 32166
rect 22008 32020 22060 32026
rect 22008 31962 22060 31968
rect 22112 31958 22140 32914
rect 22296 32570 22324 33390
rect 22284 32564 22336 32570
rect 22284 32506 22336 32512
rect 22848 32434 22876 33798
rect 23860 33318 23888 33798
rect 23848 33312 23900 33318
rect 23848 33254 23900 33260
rect 23860 32910 23888 33254
rect 23952 32978 23980 34478
rect 24872 34474 24900 35634
rect 25056 35154 25084 36094
rect 25136 36032 25188 36038
rect 25136 35974 25188 35980
rect 25148 35766 25176 35974
rect 25136 35760 25188 35766
rect 25136 35702 25188 35708
rect 25044 35148 25096 35154
rect 25044 35090 25096 35096
rect 26056 35148 26108 35154
rect 26056 35090 26108 35096
rect 24952 34740 25004 34746
rect 24952 34682 25004 34688
rect 24860 34468 24912 34474
rect 24860 34410 24912 34416
rect 24400 34400 24452 34406
rect 24400 34342 24452 34348
rect 24412 33998 24440 34342
rect 24872 34066 24900 34410
rect 24860 34060 24912 34066
rect 24860 34002 24912 34008
rect 24400 33992 24452 33998
rect 24400 33934 24452 33940
rect 24872 33522 24900 34002
rect 24216 33516 24268 33522
rect 24216 33458 24268 33464
rect 24860 33516 24912 33522
rect 24860 33458 24912 33464
rect 24228 33114 24256 33458
rect 24964 33318 24992 34682
rect 25056 34218 25084 35090
rect 25688 34944 25740 34950
rect 25688 34886 25740 34892
rect 25700 34610 25728 34886
rect 25688 34604 25740 34610
rect 25688 34546 25740 34552
rect 26068 34542 26096 35090
rect 26160 35018 26188 36722
rect 26436 36174 26464 37810
rect 26516 37664 26568 37670
rect 26516 37606 26568 37612
rect 26528 37194 26556 37606
rect 26516 37188 26568 37194
rect 26516 37130 26568 37136
rect 26700 37120 26752 37126
rect 26700 37062 26752 37068
rect 26712 36854 26740 37062
rect 26700 36848 26752 36854
rect 26700 36790 26752 36796
rect 27172 36378 27200 37810
rect 27724 37398 27752 38150
rect 28080 37868 28132 37874
rect 28080 37810 28132 37816
rect 28092 37670 28120 37810
rect 27988 37664 28040 37670
rect 27988 37606 28040 37612
rect 28080 37664 28132 37670
rect 28080 37606 28132 37612
rect 27712 37392 27764 37398
rect 27712 37334 27764 37340
rect 28000 37330 28028 37606
rect 28080 37460 28132 37466
rect 28080 37402 28132 37408
rect 27988 37324 28040 37330
rect 27988 37266 28040 37272
rect 28000 37194 28028 37266
rect 27988 37188 28040 37194
rect 27988 37130 28040 37136
rect 27988 36848 28040 36854
rect 27988 36790 28040 36796
rect 27252 36576 27304 36582
rect 27252 36518 27304 36524
rect 27160 36372 27212 36378
rect 27160 36314 27212 36320
rect 26424 36168 26476 36174
rect 26424 36110 26476 36116
rect 26976 36100 27028 36106
rect 26976 36042 27028 36048
rect 26516 36032 26568 36038
rect 26516 35974 26568 35980
rect 26528 35766 26556 35974
rect 26516 35760 26568 35766
rect 26516 35702 26568 35708
rect 26988 35222 27016 36042
rect 26976 35216 27028 35222
rect 26976 35158 27028 35164
rect 27264 35154 27292 36518
rect 27620 36236 27672 36242
rect 27620 36178 27672 36184
rect 27632 35290 27660 36178
rect 28000 36174 28028 36790
rect 27988 36168 28040 36174
rect 27988 36110 28040 36116
rect 28092 35698 28120 37402
rect 28552 36854 28580 38286
rect 28724 38208 28776 38214
rect 28724 38150 28776 38156
rect 28632 37664 28684 37670
rect 28632 37606 28684 37612
rect 28644 37262 28672 37606
rect 28632 37256 28684 37262
rect 28632 37198 28684 37204
rect 28540 36848 28592 36854
rect 28540 36790 28592 36796
rect 28172 36576 28224 36582
rect 28172 36518 28224 36524
rect 28080 35692 28132 35698
rect 28080 35634 28132 35640
rect 27712 35624 27764 35630
rect 27712 35566 27764 35572
rect 27620 35284 27672 35290
rect 27620 35226 27672 35232
rect 27252 35148 27304 35154
rect 27252 35090 27304 35096
rect 26700 35080 26752 35086
rect 26700 35022 26752 35028
rect 26148 35012 26200 35018
rect 26148 34954 26200 34960
rect 26056 34536 26108 34542
rect 26056 34478 26108 34484
rect 26240 34400 26292 34406
rect 26240 34342 26292 34348
rect 25056 34190 25176 34218
rect 24952 33312 25004 33318
rect 24952 33254 25004 33260
rect 24216 33108 24268 33114
rect 24216 33050 24268 33056
rect 23940 32972 23992 32978
rect 23940 32914 23992 32920
rect 23848 32904 23900 32910
rect 23848 32846 23900 32852
rect 23204 32768 23256 32774
rect 23204 32710 23256 32716
rect 22192 32428 22244 32434
rect 22192 32370 22244 32376
rect 22836 32428 22888 32434
rect 22836 32370 22888 32376
rect 22204 32026 22232 32370
rect 22284 32360 22336 32366
rect 22284 32302 22336 32308
rect 22192 32020 22244 32026
rect 22192 31962 22244 31968
rect 22100 31952 22152 31958
rect 22152 31900 22232 31906
rect 22100 31894 22232 31900
rect 22112 31878 22232 31894
rect 21456 31748 21508 31754
rect 21456 31690 21508 31696
rect 20904 31340 20956 31346
rect 20904 31282 20956 31288
rect 21272 31340 21324 31346
rect 21272 31282 21324 31288
rect 20812 30728 20864 30734
rect 20812 30670 20864 30676
rect 20824 30326 20852 30670
rect 20812 30320 20864 30326
rect 20916 30297 20944 31282
rect 21284 30870 21312 31282
rect 21364 31136 21416 31142
rect 21364 31078 21416 31084
rect 21272 30864 21324 30870
rect 21272 30806 21324 30812
rect 21376 30666 21404 31078
rect 22204 30802 22232 31878
rect 22192 30796 22244 30802
rect 22192 30738 22244 30744
rect 21364 30660 21416 30666
rect 21364 30602 21416 30608
rect 22296 30326 22324 32302
rect 22560 31884 22612 31890
rect 22560 31826 22612 31832
rect 22572 31754 22600 31826
rect 23216 31822 23244 32710
rect 23388 32564 23440 32570
rect 23388 32506 23440 32512
rect 23296 32224 23348 32230
rect 23296 32166 23348 32172
rect 23204 31816 23256 31822
rect 23204 31758 23256 31764
rect 22572 31726 22692 31754
rect 22664 31278 22692 31726
rect 23308 31482 23336 32166
rect 23400 31958 23428 32506
rect 23952 32366 23980 32914
rect 24964 32774 24992 33254
rect 25148 32978 25176 34190
rect 26252 34066 26280 34342
rect 26712 34202 26740 35022
rect 27264 34610 27292 35090
rect 27252 34604 27304 34610
rect 27252 34546 27304 34552
rect 27724 34202 27752 35566
rect 27896 35080 27948 35086
rect 27896 35022 27948 35028
rect 27908 34406 27936 35022
rect 28092 34762 28120 35634
rect 28184 35290 28212 36518
rect 28448 36100 28500 36106
rect 28448 36042 28500 36048
rect 28264 36032 28316 36038
rect 28264 35974 28316 35980
rect 28172 35284 28224 35290
rect 28172 35226 28224 35232
rect 28000 34734 28120 34762
rect 27896 34400 27948 34406
rect 27896 34342 27948 34348
rect 26700 34196 26752 34202
rect 26700 34138 26752 34144
rect 27712 34196 27764 34202
rect 27712 34138 27764 34144
rect 26240 34060 26292 34066
rect 26240 34002 26292 34008
rect 26608 33924 26660 33930
rect 26608 33866 26660 33872
rect 26240 33516 26292 33522
rect 26240 33458 26292 33464
rect 26252 33114 26280 33458
rect 26620 33114 26648 33866
rect 26712 33386 26740 34138
rect 27712 33448 27764 33454
rect 27712 33390 27764 33396
rect 26700 33380 26752 33386
rect 26700 33322 26752 33328
rect 26240 33108 26292 33114
rect 26240 33050 26292 33056
rect 26608 33108 26660 33114
rect 26608 33050 26660 33056
rect 26712 32978 26740 33322
rect 27528 33312 27580 33318
rect 27528 33254 27580 33260
rect 25136 32972 25188 32978
rect 25136 32914 25188 32920
rect 26700 32972 26752 32978
rect 26700 32914 26752 32920
rect 24952 32768 25004 32774
rect 24952 32710 25004 32716
rect 25148 32502 25176 32914
rect 26608 32904 26660 32910
rect 26608 32846 26660 32852
rect 25320 32836 25372 32842
rect 25320 32778 25372 32784
rect 25136 32496 25188 32502
rect 25136 32438 25188 32444
rect 23940 32360 23992 32366
rect 23940 32302 23992 32308
rect 23388 31952 23440 31958
rect 23388 31894 23440 31900
rect 23400 31822 23428 31894
rect 23388 31816 23440 31822
rect 23388 31758 23440 31764
rect 23952 31754 23980 32302
rect 25044 32292 25096 32298
rect 25044 32234 25096 32240
rect 24952 32224 25004 32230
rect 24952 32166 25004 32172
rect 24964 31890 24992 32166
rect 24952 31884 25004 31890
rect 24952 31826 25004 31832
rect 24676 31816 24728 31822
rect 24676 31758 24728 31764
rect 23952 31726 24072 31754
rect 23296 31476 23348 31482
rect 23296 31418 23348 31424
rect 23848 31340 23900 31346
rect 23848 31282 23900 31288
rect 22652 31272 22704 31278
rect 22652 31214 22704 31220
rect 22928 31272 22980 31278
rect 22928 31214 22980 31220
rect 22284 30320 22336 30326
rect 20812 30262 20864 30268
rect 20902 30288 20958 30297
rect 20824 30190 20852 30262
rect 22284 30262 22336 30268
rect 20902 30223 20958 30232
rect 22376 30252 22428 30258
rect 20812 30184 20864 30190
rect 20812 30126 20864 30132
rect 20812 28484 20864 28490
rect 20812 28426 20864 28432
rect 20824 28218 20852 28426
rect 20812 28212 20864 28218
rect 20812 28154 20864 28160
rect 20812 27600 20864 27606
rect 20812 27542 20864 27548
rect 20720 26988 20772 26994
rect 20720 26930 20772 26936
rect 20628 26444 20680 26450
rect 20824 26432 20852 27542
rect 20680 26404 20852 26432
rect 20628 26386 20680 26392
rect 20548 26302 20668 26330
rect 20640 26296 20668 26302
rect 20640 26268 20760 26296
rect 20168 25356 20220 25362
rect 20168 25298 20220 25304
rect 20180 23526 20208 25298
rect 20732 25294 20760 26268
rect 20720 25288 20772 25294
rect 20720 25230 20772 25236
rect 20352 24812 20404 24818
rect 20352 24754 20404 24760
rect 20364 24410 20392 24754
rect 20352 24404 20404 24410
rect 20352 24346 20404 24352
rect 20732 24206 20760 25230
rect 20824 24750 20852 26404
rect 20812 24744 20864 24750
rect 20812 24686 20864 24692
rect 20916 24290 20944 30223
rect 22376 30194 22428 30200
rect 21180 30048 21232 30054
rect 21180 29990 21232 29996
rect 21192 29578 21220 29990
rect 22388 29850 22416 30194
rect 22284 29844 22336 29850
rect 22284 29786 22336 29792
rect 22376 29844 22428 29850
rect 22376 29786 22428 29792
rect 21180 29572 21232 29578
rect 21180 29514 21232 29520
rect 21640 29572 21692 29578
rect 21640 29514 21692 29520
rect 21652 29306 21680 29514
rect 21640 29300 21692 29306
rect 21640 29242 21692 29248
rect 22192 29164 22244 29170
rect 22192 29106 22244 29112
rect 21272 29096 21324 29102
rect 21272 29038 21324 29044
rect 21284 27470 21312 29038
rect 22100 28960 22152 28966
rect 22100 28902 22152 28908
rect 22112 28082 22140 28902
rect 22204 28082 22232 29106
rect 22296 28150 22324 29786
rect 22664 29034 22692 31214
rect 22940 30734 22968 31214
rect 23572 31136 23624 31142
rect 23572 31078 23624 31084
rect 23584 30734 23612 31078
rect 23860 30938 23888 31282
rect 23848 30932 23900 30938
rect 23848 30874 23900 30880
rect 22928 30728 22980 30734
rect 22928 30670 22980 30676
rect 23572 30728 23624 30734
rect 23572 30670 23624 30676
rect 22940 29714 22968 30670
rect 23860 30666 23888 30874
rect 23848 30660 23900 30666
rect 23848 30602 23900 30608
rect 23860 30258 23888 30602
rect 23848 30252 23900 30258
rect 23848 30194 23900 30200
rect 24044 30190 24072 31726
rect 24584 31340 24636 31346
rect 24584 31282 24636 31288
rect 24596 30938 24624 31282
rect 24688 31278 24716 31758
rect 25056 31482 25084 32234
rect 25044 31476 25096 31482
rect 25044 31418 25096 31424
rect 24676 31272 24728 31278
rect 24676 31214 24728 31220
rect 25056 30954 25084 31418
rect 24584 30932 24636 30938
rect 24584 30874 24636 30880
rect 24964 30926 25084 30954
rect 24860 30796 24912 30802
rect 24860 30738 24912 30744
rect 24872 30190 24900 30738
rect 24964 30734 24992 30926
rect 25148 30802 25176 32438
rect 25332 32366 25360 32778
rect 26620 32434 26648 32846
rect 27540 32502 27568 33254
rect 27724 33046 27752 33390
rect 27712 33040 27764 33046
rect 27712 32982 27764 32988
rect 27528 32496 27580 32502
rect 27528 32438 27580 32444
rect 27724 32434 27752 32982
rect 28000 32910 28028 34734
rect 28184 33998 28212 35226
rect 28276 35154 28304 35974
rect 28460 35766 28488 36042
rect 28540 36032 28592 36038
rect 28540 35974 28592 35980
rect 28448 35760 28500 35766
rect 28448 35702 28500 35708
rect 28356 35488 28408 35494
rect 28356 35430 28408 35436
rect 28264 35148 28316 35154
rect 28264 35090 28316 35096
rect 28264 34944 28316 34950
rect 28264 34886 28316 34892
rect 28276 34746 28304 34886
rect 28264 34740 28316 34746
rect 28264 34682 28316 34688
rect 28276 34134 28304 34682
rect 28264 34128 28316 34134
rect 28264 34070 28316 34076
rect 28172 33992 28224 33998
rect 28172 33934 28224 33940
rect 28368 32978 28396 35430
rect 28460 35086 28488 35702
rect 28552 35290 28580 35974
rect 28632 35556 28684 35562
rect 28632 35498 28684 35504
rect 28540 35284 28592 35290
rect 28540 35226 28592 35232
rect 28448 35080 28500 35086
rect 28448 35022 28500 35028
rect 28540 35012 28592 35018
rect 28540 34954 28592 34960
rect 28448 34944 28500 34950
rect 28448 34886 28500 34892
rect 28460 34678 28488 34886
rect 28448 34672 28500 34678
rect 28448 34614 28500 34620
rect 28460 33930 28488 34614
rect 28552 33998 28580 34954
rect 28644 34746 28672 35498
rect 28632 34740 28684 34746
rect 28632 34682 28684 34688
rect 28632 34400 28684 34406
rect 28632 34342 28684 34348
rect 28644 33998 28672 34342
rect 28540 33992 28592 33998
rect 28540 33934 28592 33940
rect 28632 33992 28684 33998
rect 28632 33934 28684 33940
rect 28448 33924 28500 33930
rect 28448 33866 28500 33872
rect 28540 33856 28592 33862
rect 28540 33798 28592 33804
rect 28356 32972 28408 32978
rect 28356 32914 28408 32920
rect 27988 32904 28040 32910
rect 27988 32846 28040 32852
rect 28264 32768 28316 32774
rect 28264 32710 28316 32716
rect 26608 32428 26660 32434
rect 26608 32370 26660 32376
rect 27712 32428 27764 32434
rect 27712 32370 27764 32376
rect 25320 32360 25372 32366
rect 25320 32302 25372 32308
rect 25332 31890 25360 32302
rect 26424 32224 26476 32230
rect 26424 32166 26476 32172
rect 25320 31884 25372 31890
rect 25320 31826 25372 31832
rect 26436 31414 26464 32166
rect 26620 31754 26648 32370
rect 27712 32224 27764 32230
rect 27712 32166 27764 32172
rect 27620 31816 27672 31822
rect 27620 31758 27672 31764
rect 26608 31748 26660 31754
rect 26608 31690 26660 31696
rect 26424 31408 26476 31414
rect 26424 31350 26476 31356
rect 25136 30796 25188 30802
rect 25136 30738 25188 30744
rect 26620 30734 26648 31690
rect 26884 31680 26936 31686
rect 26884 31622 26936 31628
rect 26896 31414 26924 31622
rect 26884 31408 26936 31414
rect 26884 31350 26936 31356
rect 27632 31210 27660 31758
rect 27620 31204 27672 31210
rect 27620 31146 27672 31152
rect 24952 30728 25004 30734
rect 24952 30670 25004 30676
rect 25964 30728 26016 30734
rect 25964 30670 26016 30676
rect 26608 30728 26660 30734
rect 26608 30670 26660 30676
rect 27344 30728 27396 30734
rect 27344 30670 27396 30676
rect 27620 30728 27672 30734
rect 27620 30670 27672 30676
rect 25228 30592 25280 30598
rect 25228 30534 25280 30540
rect 25044 30252 25096 30258
rect 25044 30194 25096 30200
rect 23756 30184 23808 30190
rect 23756 30126 23808 30132
rect 24032 30184 24084 30190
rect 24032 30126 24084 30132
rect 24860 30184 24912 30190
rect 24860 30126 24912 30132
rect 23572 30116 23624 30122
rect 23572 30058 23624 30064
rect 23480 30048 23532 30054
rect 23480 29990 23532 29996
rect 22928 29708 22980 29714
rect 22928 29650 22980 29656
rect 23492 29646 23520 29990
rect 23584 29714 23612 30058
rect 23572 29708 23624 29714
rect 23572 29650 23624 29656
rect 23664 29708 23716 29714
rect 23664 29650 23716 29656
rect 23480 29640 23532 29646
rect 23480 29582 23532 29588
rect 23584 29170 23612 29650
rect 23572 29164 23624 29170
rect 23572 29106 23624 29112
rect 22836 29096 22888 29102
rect 23676 29050 23704 29650
rect 23768 29306 23796 30126
rect 23756 29300 23808 29306
rect 23756 29242 23808 29248
rect 24044 29220 24072 30126
rect 24872 30054 24900 30126
rect 24860 30048 24912 30054
rect 24860 29990 24912 29996
rect 24872 29730 24900 29990
rect 25056 29850 25084 30194
rect 25044 29844 25096 29850
rect 25044 29786 25096 29792
rect 24872 29702 24992 29730
rect 25240 29714 25268 30534
rect 25976 30394 26004 30670
rect 26516 30592 26568 30598
rect 26516 30534 26568 30540
rect 25964 30388 26016 30394
rect 25964 30330 26016 30336
rect 24860 29640 24912 29646
rect 24860 29582 24912 29588
rect 24044 29192 24164 29220
rect 24136 29102 24164 29192
rect 24872 29102 24900 29582
rect 22836 29038 22888 29044
rect 22652 29028 22704 29034
rect 22652 28970 22704 28976
rect 22848 28558 22876 29038
rect 23584 29034 23704 29050
rect 24124 29096 24176 29102
rect 24124 29038 24176 29044
rect 24860 29096 24912 29102
rect 24860 29038 24912 29044
rect 23572 29028 23704 29034
rect 23624 29022 23704 29028
rect 23572 28970 23624 28976
rect 22836 28552 22888 28558
rect 22836 28494 22888 28500
rect 23480 28484 23532 28490
rect 23480 28426 23532 28432
rect 23204 28416 23256 28422
rect 23204 28358 23256 28364
rect 22284 28144 22336 28150
rect 22284 28086 22336 28092
rect 22100 28076 22152 28082
rect 22100 28018 22152 28024
rect 22192 28076 22244 28082
rect 22192 28018 22244 28024
rect 23020 28076 23072 28082
rect 23020 28018 23072 28024
rect 22100 27872 22152 27878
rect 22100 27814 22152 27820
rect 21272 27464 21324 27470
rect 21272 27406 21324 27412
rect 21364 27328 21416 27334
rect 21364 27270 21416 27276
rect 21376 27130 21404 27270
rect 21364 27124 21416 27130
rect 21364 27066 21416 27072
rect 20996 26784 21048 26790
rect 20996 26726 21048 26732
rect 21008 26314 21036 26726
rect 22112 26382 22140 27814
rect 22204 27674 22232 28018
rect 22192 27668 22244 27674
rect 22192 27610 22244 27616
rect 22192 27328 22244 27334
rect 22192 27270 22244 27276
rect 22652 27328 22704 27334
rect 22652 27270 22704 27276
rect 22204 26994 22232 27270
rect 22664 27130 22692 27270
rect 22652 27124 22704 27130
rect 22652 27066 22704 27072
rect 22192 26988 22244 26994
rect 22192 26930 22244 26936
rect 22376 26784 22428 26790
rect 22376 26726 22428 26732
rect 22388 26586 22416 26726
rect 22664 26586 22692 27066
rect 22376 26580 22428 26586
rect 22376 26522 22428 26528
rect 22652 26580 22704 26586
rect 22652 26522 22704 26528
rect 22100 26376 22152 26382
rect 22100 26318 22152 26324
rect 20996 26308 21048 26314
rect 20996 26250 21048 26256
rect 20996 25968 21048 25974
rect 20996 25910 21048 25916
rect 21008 25498 21036 25910
rect 21088 25696 21140 25702
rect 21088 25638 21140 25644
rect 20996 25492 21048 25498
rect 20996 25434 21048 25440
rect 21100 24954 21128 25638
rect 22284 25152 22336 25158
rect 22284 25094 22336 25100
rect 21088 24948 21140 24954
rect 21088 24890 21140 24896
rect 22296 24886 22324 25094
rect 20996 24880 21048 24886
rect 20996 24822 21048 24828
rect 22284 24880 22336 24886
rect 22284 24822 22336 24828
rect 20824 24262 20944 24290
rect 20720 24200 20772 24206
rect 20720 24142 20772 24148
rect 20824 23866 20852 24262
rect 20904 24132 20956 24138
rect 20904 24074 20956 24080
rect 20812 23860 20864 23866
rect 20812 23802 20864 23808
rect 20168 23520 20220 23526
rect 20168 23462 20220 23468
rect 20180 23186 20208 23462
rect 20260 23316 20312 23322
rect 20260 23258 20312 23264
rect 20168 23180 20220 23186
rect 20168 23122 20220 23128
rect 20272 22506 20300 23258
rect 20916 22982 20944 24074
rect 21008 23322 21036 24822
rect 21824 24744 21876 24750
rect 21824 24686 21876 24692
rect 21180 24200 21232 24206
rect 21180 24142 21232 24148
rect 21088 24064 21140 24070
rect 21088 24006 21140 24012
rect 21100 23730 21128 24006
rect 21088 23724 21140 23730
rect 21088 23666 21140 23672
rect 20996 23316 21048 23322
rect 20996 23258 21048 23264
rect 20996 23180 21048 23186
rect 20996 23122 21048 23128
rect 20904 22976 20956 22982
rect 20904 22918 20956 22924
rect 20536 22636 20588 22642
rect 20536 22578 20588 22584
rect 20260 22500 20312 22506
rect 20260 22442 20312 22448
rect 20168 22432 20220 22438
rect 20168 22374 20220 22380
rect 20180 22030 20208 22374
rect 20272 22234 20300 22442
rect 20260 22228 20312 22234
rect 20260 22170 20312 22176
rect 20168 22024 20220 22030
rect 20168 21966 20220 21972
rect 20076 21004 20128 21010
rect 20076 20946 20128 20952
rect 19892 20936 19944 20942
rect 19892 20878 19944 20884
rect 19800 20392 19852 20398
rect 19800 20334 19852 20340
rect 19708 20052 19760 20058
rect 19708 19994 19760 20000
rect 18880 18964 18932 18970
rect 18880 18906 18932 18912
rect 19432 18964 19484 18970
rect 19432 18906 19484 18912
rect 18788 18692 18840 18698
rect 18788 18634 18840 18640
rect 19444 18426 19472 18906
rect 19812 18902 19840 20334
rect 19904 19378 19932 20878
rect 19892 19372 19944 19378
rect 19892 19314 19944 19320
rect 19800 18896 19852 18902
rect 19800 18838 19852 18844
rect 19432 18420 19484 18426
rect 19432 18362 19484 18368
rect 19444 17746 19472 18362
rect 19432 17740 19484 17746
rect 19432 17682 19484 17688
rect 18696 17672 18748 17678
rect 18696 17614 18748 17620
rect 18604 17604 18656 17610
rect 18604 17546 18656 17552
rect 18616 16794 18644 17546
rect 18708 17134 18736 17614
rect 18880 17536 18932 17542
rect 18880 17478 18932 17484
rect 18892 17338 18920 17478
rect 18880 17332 18932 17338
rect 20088 17320 20116 20946
rect 20272 19310 20300 22170
rect 20548 21690 20576 22578
rect 20536 21684 20588 21690
rect 20536 21626 20588 21632
rect 21008 21486 21036 23122
rect 21192 22642 21220 24142
rect 21456 23520 21508 23526
rect 21456 23462 21508 23468
rect 21468 23118 21496 23462
rect 21836 23186 21864 24686
rect 22744 24608 22796 24614
rect 22744 24550 22796 24556
rect 22560 24064 22612 24070
rect 22560 24006 22612 24012
rect 21824 23180 21876 23186
rect 21824 23122 21876 23128
rect 21456 23112 21508 23118
rect 21456 23054 21508 23060
rect 21180 22636 21232 22642
rect 21180 22578 21232 22584
rect 21088 21548 21140 21554
rect 21088 21490 21140 21496
rect 20996 21480 21048 21486
rect 20996 21422 21048 21428
rect 20720 21004 20772 21010
rect 20720 20946 20772 20952
rect 20628 20460 20680 20466
rect 20628 20402 20680 20408
rect 20640 19514 20668 20402
rect 20732 20398 20760 20946
rect 20720 20392 20772 20398
rect 20720 20334 20772 20340
rect 20720 20256 20772 20262
rect 20720 20198 20772 20204
rect 20732 19786 20760 20198
rect 20720 19780 20772 19786
rect 20720 19722 20772 19728
rect 20628 19508 20680 19514
rect 20628 19450 20680 19456
rect 20812 19508 20864 19514
rect 20812 19450 20864 19456
rect 20260 19304 20312 19310
rect 20260 19246 20312 19252
rect 20272 18834 20300 19246
rect 20260 18828 20312 18834
rect 20260 18770 20312 18776
rect 20272 18222 20300 18770
rect 20824 18426 20852 19450
rect 20904 18692 20956 18698
rect 20904 18634 20956 18640
rect 20812 18420 20864 18426
rect 20812 18362 20864 18368
rect 20916 18358 20944 18634
rect 20904 18352 20956 18358
rect 20904 18294 20956 18300
rect 20720 18284 20772 18290
rect 20720 18226 20772 18232
rect 20260 18216 20312 18222
rect 20260 18158 20312 18164
rect 20352 18080 20404 18086
rect 20352 18022 20404 18028
rect 20364 17678 20392 18022
rect 20352 17672 20404 17678
rect 20352 17614 20404 17620
rect 18880 17274 18932 17280
rect 19996 17292 20116 17320
rect 18696 17128 18748 17134
rect 18696 17070 18748 17076
rect 18880 16992 18932 16998
rect 18880 16934 18932 16940
rect 18604 16788 18656 16794
rect 18604 16730 18656 16736
rect 18892 16114 18920 16934
rect 19340 16516 19392 16522
rect 19340 16458 19392 16464
rect 19352 16250 19380 16458
rect 19340 16244 19392 16250
rect 19340 16186 19392 16192
rect 18880 16108 18932 16114
rect 18880 16050 18932 16056
rect 17408 15496 17460 15502
rect 17408 15438 17460 15444
rect 18512 15496 18564 15502
rect 18512 15438 18564 15444
rect 16304 15088 16356 15094
rect 16304 15030 16356 15036
rect 15844 14952 15896 14958
rect 15844 14894 15896 14900
rect 14740 11756 14792 11762
rect 14740 11698 14792 11704
rect 14464 11144 14516 11150
rect 14464 11086 14516 11092
rect 17224 11144 17276 11150
rect 17224 11086 17276 11092
rect 15476 10124 15528 10130
rect 15476 10066 15528 10072
rect 14280 9580 14332 9586
rect 14280 9522 14332 9528
rect 14188 9104 14240 9110
rect 14188 9046 14240 9052
rect 13912 9036 13964 9042
rect 13912 8978 13964 8984
rect 13544 8968 13596 8974
rect 13544 8910 13596 8916
rect 13636 8968 13688 8974
rect 13636 8910 13688 8916
rect 12716 8900 12768 8906
rect 12716 8842 12768 8848
rect 13556 8566 13584 8910
rect 13544 8560 13596 8566
rect 13544 8502 13596 8508
rect 13556 7886 13584 8502
rect 13648 8430 13676 8910
rect 13636 8424 13688 8430
rect 13636 8366 13688 8372
rect 13648 7954 13676 8366
rect 14200 8362 14228 9046
rect 14292 8566 14320 9522
rect 15108 9512 15160 9518
rect 15108 9454 15160 9460
rect 14556 8900 14608 8906
rect 14556 8842 14608 8848
rect 14568 8634 14596 8842
rect 14556 8628 14608 8634
rect 14556 8570 14608 8576
rect 14280 8560 14332 8566
rect 14280 8502 14332 8508
rect 14464 8492 14516 8498
rect 14464 8434 14516 8440
rect 14188 8356 14240 8362
rect 14188 8298 14240 8304
rect 14476 8090 14504 8434
rect 14556 8356 14608 8362
rect 14556 8298 14608 8304
rect 14464 8084 14516 8090
rect 14464 8026 14516 8032
rect 13636 7948 13688 7954
rect 13636 7890 13688 7896
rect 13544 7880 13596 7886
rect 13544 7822 13596 7828
rect 12624 7812 12676 7818
rect 12624 7754 12676 7760
rect 14372 7744 14424 7750
rect 14372 7686 14424 7692
rect 14384 7478 14412 7686
rect 14372 7472 14424 7478
rect 14372 7414 14424 7420
rect 9220 7404 9272 7410
rect 9220 7346 9272 7352
rect 11796 7404 11848 7410
rect 11796 7346 11848 7352
rect 12348 7404 12400 7410
rect 12348 7346 12400 7352
rect 12440 7404 12492 7410
rect 12440 7346 12492 7352
rect 11808 6798 11836 7346
rect 12164 7200 12216 7206
rect 12164 7142 12216 7148
rect 12176 7002 12204 7142
rect 12164 6996 12216 7002
rect 12164 6938 12216 6944
rect 11336 6792 11388 6798
rect 11336 6734 11388 6740
rect 11796 6792 11848 6798
rect 11796 6734 11848 6740
rect 11348 5710 11376 6734
rect 12360 6458 12388 7346
rect 12808 7200 12860 7206
rect 12808 7142 12860 7148
rect 12820 6730 12848 7142
rect 14568 6914 14596 8298
rect 15120 8106 15148 9454
rect 15488 8838 15516 10066
rect 15476 8832 15528 8838
rect 15476 8774 15528 8780
rect 16028 8832 16080 8838
rect 16028 8774 16080 8780
rect 15488 8430 15516 8774
rect 15568 8628 15620 8634
rect 15568 8570 15620 8576
rect 15476 8424 15528 8430
rect 15476 8366 15528 8372
rect 15120 8078 15240 8106
rect 15212 8022 15240 8078
rect 15200 8016 15252 8022
rect 15200 7958 15252 7964
rect 15384 8016 15436 8022
rect 15384 7958 15436 7964
rect 15292 7336 15344 7342
rect 15292 7278 15344 7284
rect 14476 6886 14596 6914
rect 12808 6724 12860 6730
rect 12808 6666 12860 6672
rect 12348 6452 12400 6458
rect 12348 6394 12400 6400
rect 11980 6316 12032 6322
rect 11980 6258 12032 6264
rect 12992 6316 13044 6322
rect 12992 6258 13044 6264
rect 11612 6112 11664 6118
rect 11612 6054 11664 6060
rect 11624 5778 11652 6054
rect 11612 5772 11664 5778
rect 11612 5714 11664 5720
rect 11336 5704 11388 5710
rect 11336 5646 11388 5652
rect 10876 5024 10928 5030
rect 10876 4966 10928 4972
rect 10784 4480 10836 4486
rect 10784 4422 10836 4428
rect 9864 3936 9916 3942
rect 9864 3878 9916 3884
rect 9876 3534 9904 3878
rect 9864 3528 9916 3534
rect 9864 3470 9916 3476
rect 10796 3466 10824 4422
rect 10888 3466 10916 4966
rect 10968 4140 11020 4146
rect 10968 4082 11020 4088
rect 10784 3460 10836 3466
rect 10784 3402 10836 3408
rect 10876 3460 10928 3466
rect 10876 3402 10928 3408
rect 7840 3052 7892 3058
rect 7840 2994 7892 3000
rect 1584 2848 1636 2854
rect 1584 2790 1636 2796
rect 1400 2304 1452 2310
rect 1400 2246 1452 2252
rect 1412 800 1440 2246
rect 1596 2009 1624 2790
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 10980 2582 11008 4082
rect 11348 3602 11376 5646
rect 11992 4826 12020 6258
rect 12624 5636 12676 5642
rect 12624 5578 12676 5584
rect 12636 5370 12664 5578
rect 13004 5370 13032 6258
rect 14476 6254 14504 6886
rect 15304 6866 15332 7278
rect 15292 6860 15344 6866
rect 15292 6802 15344 6808
rect 14740 6656 14792 6662
rect 14740 6598 14792 6604
rect 14752 6458 14780 6598
rect 14740 6452 14792 6458
rect 14740 6394 14792 6400
rect 13268 6248 13320 6254
rect 13268 6190 13320 6196
rect 14464 6248 14516 6254
rect 14464 6190 14516 6196
rect 13084 5568 13136 5574
rect 13084 5510 13136 5516
rect 12624 5364 12676 5370
rect 12624 5306 12676 5312
rect 12992 5364 13044 5370
rect 12992 5306 13044 5312
rect 13096 5234 13124 5510
rect 12624 5228 12676 5234
rect 12624 5170 12676 5176
rect 13084 5228 13136 5234
rect 13084 5170 13136 5176
rect 12072 5024 12124 5030
rect 12072 4966 12124 4972
rect 11980 4820 12032 4826
rect 11980 4762 12032 4768
rect 11888 3664 11940 3670
rect 11888 3606 11940 3612
rect 11336 3596 11388 3602
rect 11336 3538 11388 3544
rect 10968 2576 11020 2582
rect 10968 2518 11020 2524
rect 1768 2440 1820 2446
rect 1768 2382 1820 2388
rect 4436 2440 4488 2446
rect 4436 2382 4488 2388
rect 7196 2440 7248 2446
rect 7196 2382 7248 2388
rect 11152 2440 11204 2446
rect 11152 2382 11204 2388
rect 1780 2106 1808 2382
rect 4160 2304 4212 2310
rect 4160 2246 4212 2252
rect 1768 2100 1820 2106
rect 1768 2042 1820 2048
rect 1582 2000 1638 2009
rect 1582 1935 1638 1944
rect 4172 800 4200 2246
rect 4448 1970 4476 2382
rect 6920 2304 6972 2310
rect 6920 2246 6972 2252
rect 4874 2204 5182 2213
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
rect 4436 1964 4488 1970
rect 4436 1906 4488 1912
rect 6932 800 6960 2246
rect 7208 2038 7236 2382
rect 9680 2304 9732 2310
rect 9680 2246 9732 2252
rect 7196 2032 7248 2038
rect 7196 1974 7248 1980
rect 9692 800 9720 2246
rect 11164 1902 11192 2382
rect 11900 2310 11928 3606
rect 12084 3534 12112 4966
rect 12636 4486 12664 5170
rect 12716 5160 12768 5166
rect 12716 5102 12768 5108
rect 12808 5160 12860 5166
rect 12808 5102 12860 5108
rect 12348 4480 12400 4486
rect 12348 4422 12400 4428
rect 12532 4480 12584 4486
rect 12532 4422 12584 4428
rect 12624 4480 12676 4486
rect 12624 4422 12676 4428
rect 12360 4162 12388 4422
rect 12544 4282 12572 4422
rect 12532 4276 12584 4282
rect 12532 4218 12584 4224
rect 12360 4146 12480 4162
rect 12360 4140 12492 4146
rect 12360 4134 12440 4140
rect 12360 3738 12388 4134
rect 12440 4082 12492 4088
rect 12636 3942 12664 4422
rect 12728 4146 12756 5102
rect 12820 4486 12848 5102
rect 13280 4690 13308 6190
rect 14004 6180 14056 6186
rect 14004 6122 14056 6128
rect 13728 5704 13780 5710
rect 13728 5646 13780 5652
rect 13636 5228 13688 5234
rect 13636 5170 13688 5176
rect 13544 5092 13596 5098
rect 13544 5034 13596 5040
rect 13268 4684 13320 4690
rect 13268 4626 13320 4632
rect 13556 4622 13584 5034
rect 13648 4826 13676 5170
rect 13740 4826 13768 5646
rect 13636 4820 13688 4826
rect 13636 4762 13688 4768
rect 13728 4820 13780 4826
rect 13728 4762 13780 4768
rect 13544 4616 13596 4622
rect 13544 4558 13596 4564
rect 12900 4548 12952 4554
rect 12900 4490 12952 4496
rect 12808 4480 12860 4486
rect 12808 4422 12860 4428
rect 12716 4140 12768 4146
rect 12716 4082 12768 4088
rect 12624 3936 12676 3942
rect 12624 3878 12676 3884
rect 12348 3732 12400 3738
rect 12348 3674 12400 3680
rect 12164 3596 12216 3602
rect 12164 3538 12216 3544
rect 12072 3528 12124 3534
rect 12072 3470 12124 3476
rect 12176 2990 12204 3538
rect 12348 3392 12400 3398
rect 12348 3334 12400 3340
rect 12360 3126 12388 3334
rect 12348 3120 12400 3126
rect 12348 3062 12400 3068
rect 12164 2984 12216 2990
rect 12164 2926 12216 2932
rect 12176 2514 12204 2926
rect 12820 2854 12848 4422
rect 12912 4010 12940 4490
rect 13268 4072 13320 4078
rect 13268 4014 13320 4020
rect 12900 4004 12952 4010
rect 12900 3946 12952 3952
rect 12992 3936 13044 3942
rect 12992 3878 13044 3884
rect 13004 3670 13032 3878
rect 12992 3664 13044 3670
rect 12992 3606 13044 3612
rect 13280 3618 13308 4014
rect 12900 3460 12952 3466
rect 12900 3402 12952 3408
rect 12808 2848 12860 2854
rect 12808 2790 12860 2796
rect 12440 2644 12492 2650
rect 12440 2586 12492 2592
rect 12164 2508 12216 2514
rect 12164 2450 12216 2456
rect 11888 2304 11940 2310
rect 11888 2246 11940 2252
rect 11152 1896 11204 1902
rect 11152 1838 11204 1844
rect 12452 800 12480 2586
rect 12912 2378 12940 3402
rect 13004 3398 13032 3606
rect 13280 3602 13400 3618
rect 13280 3596 13412 3602
rect 13280 3590 13360 3596
rect 13360 3538 13412 3544
rect 13084 3528 13136 3534
rect 13084 3470 13136 3476
rect 12992 3392 13044 3398
rect 12992 3334 13044 3340
rect 13004 3194 13032 3334
rect 12992 3188 13044 3194
rect 12992 3130 13044 3136
rect 13096 3126 13124 3470
rect 13084 3120 13136 3126
rect 13084 3062 13136 3068
rect 13556 2514 13584 4558
rect 14016 4078 14044 6122
rect 14476 5778 14504 6190
rect 14648 6112 14700 6118
rect 14648 6054 14700 6060
rect 14464 5772 14516 5778
rect 14464 5714 14516 5720
rect 14660 5710 14688 6054
rect 14648 5704 14700 5710
rect 14648 5646 14700 5652
rect 14752 4690 14780 6394
rect 15304 5778 15332 6802
rect 15396 6390 15424 7958
rect 15488 7834 15516 8366
rect 15580 7954 15608 8570
rect 16040 8566 16068 8774
rect 16028 8560 16080 8566
rect 16028 8502 16080 8508
rect 16028 8424 16080 8430
rect 16028 8366 16080 8372
rect 17132 8424 17184 8430
rect 17132 8366 17184 8372
rect 15568 7948 15620 7954
rect 15568 7890 15620 7896
rect 15488 7806 15608 7834
rect 15476 7744 15528 7750
rect 15476 7686 15528 7692
rect 15488 7206 15516 7686
rect 15476 7200 15528 7206
rect 15476 7142 15528 7148
rect 15384 6384 15436 6390
rect 15384 6326 15436 6332
rect 15384 6248 15436 6254
rect 15384 6190 15436 6196
rect 15292 5772 15344 5778
rect 15292 5714 15344 5720
rect 15292 5636 15344 5642
rect 15292 5578 15344 5584
rect 15304 5302 15332 5578
rect 15292 5296 15344 5302
rect 15292 5238 15344 5244
rect 15396 4690 15424 6190
rect 15488 5846 15516 7142
rect 15580 6254 15608 7806
rect 15936 7404 15988 7410
rect 15936 7346 15988 7352
rect 15568 6248 15620 6254
rect 15568 6190 15620 6196
rect 15752 6248 15804 6254
rect 15752 6190 15804 6196
rect 15764 5846 15792 6190
rect 15948 5914 15976 7346
rect 16040 7342 16068 8366
rect 16304 8288 16356 8294
rect 16304 8230 16356 8236
rect 16316 7886 16344 8230
rect 17144 8090 17172 8366
rect 17132 8084 17184 8090
rect 17132 8026 17184 8032
rect 17236 7886 17264 11086
rect 16304 7880 16356 7886
rect 16304 7822 16356 7828
rect 17224 7880 17276 7886
rect 17224 7822 17276 7828
rect 16212 7812 16264 7818
rect 16212 7754 16264 7760
rect 16028 7336 16080 7342
rect 16028 7278 16080 7284
rect 16224 6798 16252 7754
rect 16212 6792 16264 6798
rect 16212 6734 16264 6740
rect 16856 6792 16908 6798
rect 16856 6734 16908 6740
rect 16120 6656 16172 6662
rect 16120 6598 16172 6604
rect 15936 5908 15988 5914
rect 15936 5850 15988 5856
rect 15476 5840 15528 5846
rect 15476 5782 15528 5788
rect 15752 5840 15804 5846
rect 15752 5782 15804 5788
rect 16132 5778 16160 6598
rect 16868 6458 16896 6734
rect 16856 6452 16908 6458
rect 16856 6394 16908 6400
rect 17236 6304 17264 7822
rect 17316 6316 17368 6322
rect 17236 6276 17316 6304
rect 17316 6258 17368 6264
rect 16856 6112 16908 6118
rect 16856 6054 16908 6060
rect 15568 5772 15620 5778
rect 15568 5714 15620 5720
rect 16120 5772 16172 5778
rect 16120 5714 16172 5720
rect 15580 5234 15608 5714
rect 16868 5642 16896 6054
rect 16856 5636 16908 5642
rect 16856 5578 16908 5584
rect 15568 5228 15620 5234
rect 15568 5170 15620 5176
rect 17040 5228 17092 5234
rect 17040 5170 17092 5176
rect 15476 5024 15528 5030
rect 15476 4966 15528 4972
rect 14740 4684 14792 4690
rect 14740 4626 14792 4632
rect 14832 4684 14884 4690
rect 14832 4626 14884 4632
rect 15384 4684 15436 4690
rect 15384 4626 15436 4632
rect 14556 4548 14608 4554
rect 14556 4490 14608 4496
rect 14568 4214 14596 4490
rect 14556 4208 14608 4214
rect 14556 4150 14608 4156
rect 14568 4078 14596 4150
rect 14004 4072 14056 4078
rect 14004 4014 14056 4020
rect 14556 4072 14608 4078
rect 14556 4014 14608 4020
rect 14016 3670 14044 4014
rect 14004 3664 14056 3670
rect 14004 3606 14056 3612
rect 14568 3534 14596 4014
rect 14844 3602 14872 4626
rect 15488 4214 15516 4966
rect 15580 4298 15608 5170
rect 16856 5024 16908 5030
rect 16856 4966 16908 4972
rect 15936 4480 15988 4486
rect 15936 4422 15988 4428
rect 16212 4480 16264 4486
rect 16212 4422 16264 4428
rect 15580 4282 15700 4298
rect 15580 4276 15712 4282
rect 15580 4270 15660 4276
rect 15660 4218 15712 4224
rect 15476 4208 15528 4214
rect 15476 4150 15528 4156
rect 14832 3596 14884 3602
rect 14832 3538 14884 3544
rect 14556 3528 14608 3534
rect 14556 3470 14608 3476
rect 14556 3392 14608 3398
rect 14556 3334 14608 3340
rect 14568 2854 14596 3334
rect 14924 3052 14976 3058
rect 14924 2994 14976 3000
rect 14556 2848 14608 2854
rect 14556 2790 14608 2796
rect 13544 2508 13596 2514
rect 13544 2450 13596 2456
rect 12900 2372 12952 2378
rect 12900 2314 12952 2320
rect 13556 1902 13584 2450
rect 14568 2038 14596 2790
rect 14936 2650 14964 2994
rect 15292 2984 15344 2990
rect 15292 2926 15344 2932
rect 14924 2644 14976 2650
rect 14924 2586 14976 2592
rect 14556 2032 14608 2038
rect 14556 1974 14608 1980
rect 13544 1896 13596 1902
rect 13544 1838 13596 1844
rect 15304 1442 15332 2926
rect 15948 2446 15976 4422
rect 16028 4072 16080 4078
rect 16028 4014 16080 4020
rect 16040 2650 16068 4014
rect 16224 3738 16252 4422
rect 16304 4140 16356 4146
rect 16304 4082 16356 4088
rect 16212 3732 16264 3738
rect 16212 3674 16264 3680
rect 16316 3058 16344 4082
rect 16868 3126 16896 4966
rect 17052 3670 17080 5170
rect 17328 4554 17356 6258
rect 17420 4690 17448 15438
rect 19996 15094 20024 17292
rect 20444 17264 20496 17270
rect 20444 17206 20496 17212
rect 20168 16516 20220 16522
rect 20168 16458 20220 16464
rect 20180 16250 20208 16458
rect 20456 16250 20484 17206
rect 20732 17134 20760 18226
rect 21008 18222 21036 21422
rect 21100 19446 21128 21490
rect 21192 20466 21220 22578
rect 21836 21486 21864 23122
rect 22572 23050 22600 24006
rect 22652 23180 22704 23186
rect 22756 23168 22784 24550
rect 23032 23746 23060 28018
rect 23216 27470 23244 28358
rect 23492 27606 23520 28426
rect 23480 27600 23532 27606
rect 23480 27542 23532 27548
rect 23204 27464 23256 27470
rect 23204 27406 23256 27412
rect 23480 27464 23532 27470
rect 23584 27418 23612 28970
rect 24136 28626 24164 29038
rect 24124 28620 24176 28626
rect 24124 28562 24176 28568
rect 24136 28014 24164 28562
rect 24584 28416 24636 28422
rect 24584 28358 24636 28364
rect 24216 28076 24268 28082
rect 24216 28018 24268 28024
rect 24124 28008 24176 28014
rect 24124 27950 24176 27956
rect 23848 27872 23900 27878
rect 23848 27814 23900 27820
rect 23664 27532 23716 27538
rect 23664 27474 23716 27480
rect 23532 27412 23612 27418
rect 23480 27406 23612 27412
rect 23492 27390 23612 27406
rect 23492 26450 23520 27390
rect 23676 27062 23704 27474
rect 23664 27056 23716 27062
rect 23664 26998 23716 27004
rect 23676 26518 23704 26998
rect 23664 26512 23716 26518
rect 23664 26454 23716 26460
rect 23480 26444 23532 26450
rect 23480 26386 23532 26392
rect 23756 26444 23808 26450
rect 23756 26386 23808 26392
rect 23480 26240 23532 26246
rect 23480 26182 23532 26188
rect 23768 26194 23796 26386
rect 23860 26382 23888 27814
rect 24228 27130 24256 28018
rect 24596 27334 24624 28358
rect 24768 28144 24820 28150
rect 24768 28086 24820 28092
rect 24676 27464 24728 27470
rect 24676 27406 24728 27412
rect 24584 27328 24636 27334
rect 24584 27270 24636 27276
rect 24216 27124 24268 27130
rect 24216 27066 24268 27072
rect 24596 27062 24624 27270
rect 24584 27056 24636 27062
rect 24584 26998 24636 27004
rect 24688 26450 24716 27406
rect 24676 26444 24728 26450
rect 24676 26386 24728 26392
rect 23848 26376 23900 26382
rect 23848 26318 23900 26324
rect 24584 26240 24636 26246
rect 23492 25770 23520 26182
rect 23768 26166 23888 26194
rect 24584 26182 24636 26188
rect 23756 26036 23808 26042
rect 23756 25978 23808 25984
rect 23480 25764 23532 25770
rect 23480 25706 23532 25712
rect 23768 25362 23796 25978
rect 23860 25362 23888 26166
rect 24596 25838 24624 26182
rect 24584 25832 24636 25838
rect 24584 25774 24636 25780
rect 24492 25696 24544 25702
rect 24492 25638 24544 25644
rect 23756 25356 23808 25362
rect 23756 25298 23808 25304
rect 23848 25356 23900 25362
rect 23848 25298 23900 25304
rect 23768 24954 23796 25298
rect 23756 24948 23808 24954
rect 23756 24890 23808 24896
rect 23664 24812 23716 24818
rect 23664 24754 23716 24760
rect 23676 24410 23704 24754
rect 23664 24404 23716 24410
rect 23664 24346 23716 24352
rect 23112 24200 23164 24206
rect 23112 24142 23164 24148
rect 23124 23866 23152 24142
rect 23112 23860 23164 23866
rect 23112 23802 23164 23808
rect 22836 23724 22888 23730
rect 23032 23718 23152 23746
rect 22836 23666 22888 23672
rect 22704 23140 22784 23168
rect 22652 23122 22704 23128
rect 22560 23044 22612 23050
rect 22560 22986 22612 22992
rect 21916 22772 21968 22778
rect 21916 22714 21968 22720
rect 21824 21480 21876 21486
rect 21824 21422 21876 21428
rect 21836 21010 21864 21422
rect 21928 21418 21956 22714
rect 22756 22642 22784 23140
rect 22744 22636 22796 22642
rect 22744 22578 22796 22584
rect 22100 22432 22152 22438
rect 22100 22374 22152 22380
rect 22112 22030 22140 22374
rect 22848 22094 22876 23666
rect 23020 22568 23072 22574
rect 23020 22510 23072 22516
rect 22664 22066 22876 22094
rect 22100 22024 22152 22030
rect 22100 21966 22152 21972
rect 22008 21888 22060 21894
rect 22008 21830 22060 21836
rect 22020 21690 22048 21830
rect 22008 21684 22060 21690
rect 22008 21626 22060 21632
rect 21916 21412 21968 21418
rect 21916 21354 21968 21360
rect 21824 21004 21876 21010
rect 21824 20946 21876 20952
rect 21364 20868 21416 20874
rect 21364 20810 21416 20816
rect 22100 20868 22152 20874
rect 22100 20810 22152 20816
rect 21180 20460 21232 20466
rect 21180 20402 21232 20408
rect 21192 20058 21220 20402
rect 21272 20256 21324 20262
rect 21272 20198 21324 20204
rect 21180 20052 21232 20058
rect 21180 19994 21232 20000
rect 21284 19786 21312 20198
rect 21272 19780 21324 19786
rect 21272 19722 21324 19728
rect 21088 19440 21140 19446
rect 21088 19382 21140 19388
rect 20996 18216 21048 18222
rect 20996 18158 21048 18164
rect 21100 17610 21128 19382
rect 21088 17604 21140 17610
rect 21088 17546 21140 17552
rect 21100 17338 21128 17546
rect 21180 17536 21232 17542
rect 21180 17478 21232 17484
rect 21088 17332 21140 17338
rect 21088 17274 21140 17280
rect 21192 17270 21220 17478
rect 21180 17264 21232 17270
rect 21180 17206 21232 17212
rect 20720 17128 20772 17134
rect 20720 17070 20772 17076
rect 20732 16794 20760 17070
rect 20720 16788 20772 16794
rect 20720 16730 20772 16736
rect 20168 16244 20220 16250
rect 20168 16186 20220 16192
rect 20444 16244 20496 16250
rect 20444 16186 20496 16192
rect 19984 15088 20036 15094
rect 19984 15030 20036 15036
rect 18696 12776 18748 12782
rect 18696 12718 18748 12724
rect 17868 11756 17920 11762
rect 17868 11698 17920 11704
rect 17880 10674 17908 11698
rect 17868 10668 17920 10674
rect 17868 10610 17920 10616
rect 18420 10600 18472 10606
rect 18420 10542 18472 10548
rect 18144 8560 18196 8566
rect 18144 8502 18196 8508
rect 18156 8090 18184 8502
rect 18144 8084 18196 8090
rect 18144 8026 18196 8032
rect 17592 6384 17644 6390
rect 17592 6326 17644 6332
rect 17604 5574 17632 6326
rect 17592 5568 17644 5574
rect 17592 5510 17644 5516
rect 17408 4684 17460 4690
rect 17408 4626 17460 4632
rect 17316 4548 17368 4554
rect 17316 4490 17368 4496
rect 17040 3664 17092 3670
rect 17040 3606 17092 3612
rect 16856 3120 16908 3126
rect 16856 3062 16908 3068
rect 16304 3052 16356 3058
rect 16304 2994 16356 3000
rect 16028 2644 16080 2650
rect 16028 2586 16080 2592
rect 17328 2446 17356 4490
rect 17500 4072 17552 4078
rect 17500 4014 17552 4020
rect 17512 3738 17540 4014
rect 17500 3732 17552 3738
rect 17500 3674 17552 3680
rect 17408 2984 17460 2990
rect 17408 2926 17460 2932
rect 17420 2650 17448 2926
rect 17408 2644 17460 2650
rect 17408 2586 17460 2592
rect 17604 2582 17632 5510
rect 18432 5234 18460 10542
rect 18420 5228 18472 5234
rect 18420 5170 18472 5176
rect 18604 5228 18656 5234
rect 18604 5170 18656 5176
rect 18144 5024 18196 5030
rect 18144 4966 18196 4972
rect 17960 4548 18012 4554
rect 17960 4490 18012 4496
rect 17972 3482 18000 4490
rect 18052 4480 18104 4486
rect 18052 4422 18104 4428
rect 18064 3534 18092 4422
rect 18156 4214 18184 4966
rect 18616 4554 18644 5170
rect 18708 4826 18736 12718
rect 18696 4820 18748 4826
rect 18696 4762 18748 4768
rect 19984 4616 20036 4622
rect 19984 4558 20036 4564
rect 18604 4548 18656 4554
rect 18604 4490 18656 4496
rect 18420 4480 18472 4486
rect 18420 4422 18472 4428
rect 18880 4480 18932 4486
rect 18880 4422 18932 4428
rect 19616 4480 19668 4486
rect 19616 4422 19668 4428
rect 18144 4208 18196 4214
rect 18144 4150 18196 4156
rect 18432 3738 18460 4422
rect 18892 4282 18920 4422
rect 18880 4276 18932 4282
rect 18880 4218 18932 4224
rect 19628 4214 19656 4422
rect 19616 4208 19668 4214
rect 19616 4150 19668 4156
rect 18420 3732 18472 3738
rect 18420 3674 18472 3680
rect 17880 3454 18000 3482
rect 18052 3528 18104 3534
rect 18052 3470 18104 3476
rect 19800 3460 19852 3466
rect 17880 3398 17908 3454
rect 19800 3402 19852 3408
rect 19892 3460 19944 3466
rect 19892 3402 19944 3408
rect 17868 3392 17920 3398
rect 17868 3334 17920 3340
rect 18604 3392 18656 3398
rect 18604 3334 18656 3340
rect 17592 2576 17644 2582
rect 17592 2518 17644 2524
rect 17880 2514 17908 3334
rect 18616 2854 18644 3334
rect 18696 3120 18748 3126
rect 18696 3062 18748 3068
rect 18052 2848 18104 2854
rect 18052 2790 18104 2796
rect 18604 2848 18656 2854
rect 18604 2790 18656 2796
rect 17868 2508 17920 2514
rect 17868 2450 17920 2456
rect 15936 2440 15988 2446
rect 15936 2382 15988 2388
rect 17316 2440 17368 2446
rect 17316 2382 17368 2388
rect 18064 2378 18092 2790
rect 18708 2650 18736 3062
rect 19812 3058 19840 3402
rect 19904 3194 19932 3402
rect 19996 3194 20024 4558
rect 20628 4480 20680 4486
rect 20628 4422 20680 4428
rect 20640 4214 20668 4422
rect 20628 4208 20680 4214
rect 20628 4150 20680 4156
rect 20628 3936 20680 3942
rect 20628 3878 20680 3884
rect 19892 3188 19944 3194
rect 19892 3130 19944 3136
rect 19984 3188 20036 3194
rect 19984 3130 20036 3136
rect 19708 3052 19760 3058
rect 19708 2994 19760 3000
rect 19800 3052 19852 3058
rect 19800 2994 19852 3000
rect 20536 3052 20588 3058
rect 20640 3040 20668 3878
rect 21376 3194 21404 20810
rect 21824 20800 21876 20806
rect 21824 20742 21876 20748
rect 21836 20534 21864 20742
rect 21824 20528 21876 20534
rect 21824 20470 21876 20476
rect 22008 20392 22060 20398
rect 22008 20334 22060 20340
rect 22020 19922 22048 20334
rect 22008 19916 22060 19922
rect 22008 19858 22060 19864
rect 22020 19378 22048 19858
rect 22008 19372 22060 19378
rect 22008 19314 22060 19320
rect 22020 18834 22048 19314
rect 22008 18828 22060 18834
rect 22008 18770 22060 18776
rect 21916 18692 21968 18698
rect 21916 18634 21968 18640
rect 21928 18426 21956 18634
rect 21916 18420 21968 18426
rect 21916 18362 21968 18368
rect 21928 17678 21956 18362
rect 22020 18222 22048 18770
rect 22112 18766 22140 20810
rect 22284 20800 22336 20806
rect 22284 20742 22336 20748
rect 22296 20058 22324 20742
rect 22560 20460 22612 20466
rect 22560 20402 22612 20408
rect 22376 20256 22428 20262
rect 22376 20198 22428 20204
rect 22284 20052 22336 20058
rect 22284 19994 22336 20000
rect 22296 19514 22324 19994
rect 22284 19508 22336 19514
rect 22284 19450 22336 19456
rect 22388 19446 22416 20198
rect 22572 20058 22600 20402
rect 22560 20052 22612 20058
rect 22560 19994 22612 20000
rect 22376 19440 22428 19446
rect 22376 19382 22428 19388
rect 22100 18760 22152 18766
rect 22100 18702 22152 18708
rect 22008 18216 22060 18222
rect 22008 18158 22060 18164
rect 22284 18216 22336 18222
rect 22284 18158 22336 18164
rect 21916 17672 21968 17678
rect 21916 17614 21968 17620
rect 21640 17128 21692 17134
rect 21640 17070 21692 17076
rect 21652 16658 21680 17070
rect 21640 16652 21692 16658
rect 21640 16594 21692 16600
rect 21652 15502 21680 16594
rect 21928 16538 21956 17614
rect 22020 17134 22048 18158
rect 22296 17882 22324 18158
rect 22284 17876 22336 17882
rect 22284 17818 22336 17824
rect 22008 17128 22060 17134
rect 22008 17070 22060 17076
rect 22284 17128 22336 17134
rect 22284 17070 22336 17076
rect 22296 16794 22324 17070
rect 22284 16788 22336 16794
rect 22284 16730 22336 16736
rect 21928 16510 22048 16538
rect 21916 15904 21968 15910
rect 21916 15846 21968 15852
rect 21928 15570 21956 15846
rect 21916 15564 21968 15570
rect 21916 15506 21968 15512
rect 21640 15496 21692 15502
rect 21640 15438 21692 15444
rect 21652 14482 21680 15438
rect 22020 15026 22048 16510
rect 22664 15570 22692 22066
rect 23032 21894 23060 22510
rect 23020 21888 23072 21894
rect 23020 21830 23072 21836
rect 22928 18624 22980 18630
rect 22928 18566 22980 18572
rect 22940 18358 22968 18566
rect 22928 18352 22980 18358
rect 22928 18294 22980 18300
rect 22744 17536 22796 17542
rect 22744 17478 22796 17484
rect 22756 17270 22784 17478
rect 22744 17264 22796 17270
rect 22744 17206 22796 17212
rect 23124 16522 23152 23718
rect 23860 23662 23888 25298
rect 24504 25294 24532 25638
rect 24492 25288 24544 25294
rect 24492 25230 24544 25236
rect 24688 25226 24716 26386
rect 24780 25906 24808 28086
rect 24872 27538 24900 29038
rect 24964 28626 24992 29702
rect 25228 29708 25280 29714
rect 25228 29650 25280 29656
rect 26528 29578 26556 30534
rect 26516 29572 26568 29578
rect 26516 29514 26568 29520
rect 26516 29232 26568 29238
rect 26516 29174 26568 29180
rect 25136 29096 25188 29102
rect 25136 29038 25188 29044
rect 25148 28762 25176 29038
rect 26528 28762 26556 29174
rect 25136 28756 25188 28762
rect 25136 28698 25188 28704
rect 26516 28756 26568 28762
rect 26516 28698 26568 28704
rect 24952 28620 25004 28626
rect 24952 28562 25004 28568
rect 25136 28620 25188 28626
rect 25136 28562 25188 28568
rect 25148 28014 25176 28562
rect 26620 28558 26648 30670
rect 27252 30660 27304 30666
rect 27252 30602 27304 30608
rect 27264 30258 27292 30602
rect 27356 30394 27384 30670
rect 27344 30388 27396 30394
rect 27344 30330 27396 30336
rect 26792 30252 26844 30258
rect 26792 30194 26844 30200
rect 27252 30252 27304 30258
rect 27252 30194 27304 30200
rect 26804 29510 26832 30194
rect 26792 29504 26844 29510
rect 26792 29446 26844 29452
rect 26700 29300 26752 29306
rect 26700 29242 26752 29248
rect 26608 28552 26660 28558
rect 26608 28494 26660 28500
rect 26620 28082 26648 28494
rect 26608 28076 26660 28082
rect 26608 28018 26660 28024
rect 25136 28008 25188 28014
rect 25136 27950 25188 27956
rect 24860 27532 24912 27538
rect 24860 27474 24912 27480
rect 24952 27396 25004 27402
rect 24952 27338 25004 27344
rect 24964 26586 24992 27338
rect 25148 26926 25176 27950
rect 26148 27872 26200 27878
rect 26148 27814 26200 27820
rect 25228 27396 25280 27402
rect 25228 27338 25280 27344
rect 25240 27130 25268 27338
rect 25228 27124 25280 27130
rect 25228 27066 25280 27072
rect 26160 26994 26188 27814
rect 26148 26988 26200 26994
rect 26148 26930 26200 26936
rect 26620 26926 26648 28018
rect 26712 26994 26740 29242
rect 26700 26988 26752 26994
rect 26700 26930 26752 26936
rect 25136 26920 25188 26926
rect 25136 26862 25188 26868
rect 26608 26920 26660 26926
rect 26608 26862 26660 26868
rect 24952 26580 25004 26586
rect 24952 26522 25004 26528
rect 26240 26444 26292 26450
rect 26240 26386 26292 26392
rect 25320 26308 25372 26314
rect 25320 26250 25372 26256
rect 25332 25974 25360 26250
rect 26056 26240 26108 26246
rect 26056 26182 26108 26188
rect 26068 26042 26096 26182
rect 26056 26036 26108 26042
rect 26056 25978 26108 25984
rect 25320 25968 25372 25974
rect 25320 25910 25372 25916
rect 24768 25900 24820 25906
rect 24768 25842 24820 25848
rect 25596 25832 25648 25838
rect 25596 25774 25648 25780
rect 24952 25696 25004 25702
rect 24952 25638 25004 25644
rect 24964 25294 24992 25638
rect 24952 25288 25004 25294
rect 24952 25230 25004 25236
rect 24676 25220 24728 25226
rect 24676 25162 24728 25168
rect 24492 25152 24544 25158
rect 24492 25094 24544 25100
rect 24860 25152 24912 25158
rect 24860 25094 24912 25100
rect 24504 24206 24532 25094
rect 24872 24954 24900 25094
rect 24860 24948 24912 24954
rect 24860 24890 24912 24896
rect 25504 24948 25556 24954
rect 25504 24890 25556 24896
rect 25516 24206 25544 24890
rect 25608 24274 25636 25774
rect 25688 25152 25740 25158
rect 25688 25094 25740 25100
rect 25872 25152 25924 25158
rect 25872 25094 25924 25100
rect 25700 24834 25728 25094
rect 25884 24886 25912 25094
rect 25872 24880 25924 24886
rect 25700 24818 25820 24834
rect 25872 24822 25924 24828
rect 25700 24812 25832 24818
rect 25700 24806 25780 24812
rect 25780 24754 25832 24760
rect 26252 24274 26280 26386
rect 26332 26240 26384 26246
rect 26332 26182 26384 26188
rect 26344 25974 26372 26182
rect 26332 25968 26384 25974
rect 26332 25910 26384 25916
rect 25596 24268 25648 24274
rect 25596 24210 25648 24216
rect 25872 24268 25924 24274
rect 25872 24210 25924 24216
rect 26240 24268 26292 24274
rect 26240 24210 26292 24216
rect 24492 24200 24544 24206
rect 24492 24142 24544 24148
rect 25504 24200 25556 24206
rect 25504 24142 25556 24148
rect 24400 24064 24452 24070
rect 24400 24006 24452 24012
rect 24412 23866 24440 24006
rect 24400 23860 24452 23866
rect 24400 23802 24452 23808
rect 23848 23656 23900 23662
rect 23848 23598 23900 23604
rect 23572 23044 23624 23050
rect 23572 22986 23624 22992
rect 23584 22098 23612 22986
rect 23664 22704 23716 22710
rect 23664 22646 23716 22652
rect 23572 22092 23624 22098
rect 23572 22034 23624 22040
rect 23572 21956 23624 21962
rect 23572 21898 23624 21904
rect 23584 21554 23612 21898
rect 23676 21690 23704 22646
rect 24504 22030 24532 24142
rect 24676 23656 24728 23662
rect 24676 23598 24728 23604
rect 24688 22642 24716 23598
rect 25608 23186 25636 24210
rect 25884 23662 25912 24210
rect 26148 24064 26200 24070
rect 26148 24006 26200 24012
rect 26160 23866 26188 24006
rect 26148 23860 26200 23866
rect 26148 23802 26200 23808
rect 25688 23656 25740 23662
rect 25688 23598 25740 23604
rect 25872 23656 25924 23662
rect 25872 23598 25924 23604
rect 26056 23656 26108 23662
rect 26056 23598 26108 23604
rect 25596 23180 25648 23186
rect 25596 23122 25648 23128
rect 25320 22976 25372 22982
rect 25320 22918 25372 22924
rect 25332 22778 25360 22918
rect 25320 22772 25372 22778
rect 25320 22714 25372 22720
rect 24676 22636 24728 22642
rect 24676 22578 24728 22584
rect 25412 22568 25464 22574
rect 25412 22510 25464 22516
rect 24952 22432 25004 22438
rect 24952 22374 25004 22380
rect 24964 22098 24992 22374
rect 24952 22092 25004 22098
rect 24952 22034 25004 22040
rect 24492 22024 24544 22030
rect 24492 21966 24544 21972
rect 23664 21684 23716 21690
rect 23664 21626 23716 21632
rect 24504 21554 24532 21966
rect 25424 21962 25452 22510
rect 25412 21956 25464 21962
rect 25412 21898 25464 21904
rect 24676 21888 24728 21894
rect 24676 21830 24728 21836
rect 23572 21548 23624 21554
rect 23572 21490 23624 21496
rect 24492 21548 24544 21554
rect 24492 21490 24544 21496
rect 23584 21010 23612 21490
rect 24308 21344 24360 21350
rect 24308 21286 24360 21292
rect 23572 21004 23624 21010
rect 23572 20946 23624 20952
rect 23756 19712 23808 19718
rect 23756 19654 23808 19660
rect 23768 19514 23796 19654
rect 23756 19508 23808 19514
rect 23756 19450 23808 19456
rect 24320 19446 24348 21286
rect 24688 20534 24716 21830
rect 25424 21690 25452 21898
rect 25412 21684 25464 21690
rect 25412 21626 25464 21632
rect 25608 21486 25636 23122
rect 25700 22098 25728 23598
rect 26068 23118 26096 23598
rect 26332 23520 26384 23526
rect 26332 23462 26384 23468
rect 26344 23118 26372 23462
rect 26056 23112 26108 23118
rect 26056 23054 26108 23060
rect 26332 23112 26384 23118
rect 26332 23054 26384 23060
rect 25964 22976 26016 22982
rect 25964 22918 26016 22924
rect 25688 22092 25740 22098
rect 25688 22034 25740 22040
rect 25596 21480 25648 21486
rect 25596 21422 25648 21428
rect 24952 21344 25004 21350
rect 24952 21286 25004 21292
rect 24964 20942 24992 21286
rect 25700 21010 25728 22034
rect 25976 22030 26004 22918
rect 26148 22636 26200 22642
rect 26148 22578 26200 22584
rect 25964 22024 26016 22030
rect 25964 21966 26016 21972
rect 26160 21894 26188 22578
rect 26712 22094 26740 26930
rect 26804 24834 26832 29446
rect 26884 29028 26936 29034
rect 26884 28970 26936 28976
rect 26896 28694 26924 28970
rect 26884 28688 26936 28694
rect 26884 28630 26936 28636
rect 26896 28490 26924 28630
rect 26884 28484 26936 28490
rect 26884 28426 26936 28432
rect 27160 27464 27212 27470
rect 27160 27406 27212 27412
rect 26884 27396 26936 27402
rect 26884 27338 26936 27344
rect 26896 26586 26924 27338
rect 26884 26580 26936 26586
rect 26884 26522 26936 26528
rect 27172 25838 27200 27406
rect 27160 25832 27212 25838
rect 27160 25774 27212 25780
rect 27172 25378 27200 25774
rect 26988 25362 27200 25378
rect 26976 25356 27200 25362
rect 27028 25350 27200 25356
rect 26976 25298 27028 25304
rect 26884 25220 26936 25226
rect 26884 25162 26936 25168
rect 26896 24954 26924 25162
rect 26884 24948 26936 24954
rect 26884 24890 26936 24896
rect 26804 24806 26924 24834
rect 26712 22066 26832 22094
rect 26148 21888 26200 21894
rect 26148 21830 26200 21836
rect 26516 21548 26568 21554
rect 26516 21490 26568 21496
rect 25780 21480 25832 21486
rect 25780 21422 25832 21428
rect 25136 21004 25188 21010
rect 25136 20946 25188 20952
rect 25320 21004 25372 21010
rect 25320 20946 25372 20952
rect 25688 21004 25740 21010
rect 25688 20946 25740 20952
rect 24952 20936 25004 20942
rect 24952 20878 25004 20884
rect 24768 20800 24820 20806
rect 24768 20742 24820 20748
rect 24676 20528 24728 20534
rect 24676 20470 24728 20476
rect 24584 20392 24636 20398
rect 24584 20334 24636 20340
rect 24596 20058 24624 20334
rect 24584 20052 24636 20058
rect 24584 19994 24636 20000
rect 24780 19854 24808 20742
rect 25148 19990 25176 20946
rect 25332 20534 25360 20946
rect 25596 20800 25648 20806
rect 25596 20742 25648 20748
rect 25608 20602 25636 20742
rect 25596 20596 25648 20602
rect 25596 20538 25648 20544
rect 25320 20528 25372 20534
rect 25320 20470 25372 20476
rect 25228 20256 25280 20262
rect 25228 20198 25280 20204
rect 25136 19984 25188 19990
rect 25136 19926 25188 19932
rect 24768 19848 24820 19854
rect 24768 19790 24820 19796
rect 25044 19712 25096 19718
rect 25044 19654 25096 19660
rect 25056 19446 25084 19654
rect 24308 19440 24360 19446
rect 24308 19382 24360 19388
rect 25044 19440 25096 19446
rect 25044 19382 25096 19388
rect 23940 19168 23992 19174
rect 23940 19110 23992 19116
rect 23952 18766 23980 19110
rect 25056 18970 25084 19382
rect 25148 19310 25176 19926
rect 25240 19922 25268 20198
rect 25332 19922 25360 20470
rect 25792 20398 25820 21422
rect 26528 21146 26556 21490
rect 26516 21140 26568 21146
rect 26516 21082 26568 21088
rect 26804 21078 26832 22066
rect 26792 21072 26844 21078
rect 26792 21014 26844 21020
rect 25780 20392 25832 20398
rect 25780 20334 25832 20340
rect 25228 19916 25280 19922
rect 25228 19858 25280 19864
rect 25320 19916 25372 19922
rect 25320 19858 25372 19864
rect 25332 19802 25360 19858
rect 25240 19774 25360 19802
rect 25136 19304 25188 19310
rect 25136 19246 25188 19252
rect 25044 18964 25096 18970
rect 25044 18906 25096 18912
rect 23940 18760 23992 18766
rect 23940 18702 23992 18708
rect 25056 18358 25084 18906
rect 25044 18352 25096 18358
rect 25044 18294 25096 18300
rect 23664 18080 23716 18086
rect 23664 18022 23716 18028
rect 24860 18080 24912 18086
rect 24860 18022 24912 18028
rect 23676 17746 23704 18022
rect 23664 17740 23716 17746
rect 23664 17682 23716 17688
rect 23388 17672 23440 17678
rect 23388 17614 23440 17620
rect 23400 16726 23428 17614
rect 23676 17338 23704 17682
rect 24872 17610 24900 18022
rect 25148 17746 25176 19246
rect 25240 17746 25268 19774
rect 25792 19242 25820 20334
rect 26424 19848 26476 19854
rect 26424 19790 26476 19796
rect 25872 19712 25924 19718
rect 25872 19654 25924 19660
rect 25884 19310 25912 19654
rect 26436 19378 26464 19790
rect 26792 19712 26844 19718
rect 26792 19654 26844 19660
rect 26424 19372 26476 19378
rect 26424 19314 26476 19320
rect 25872 19304 25924 19310
rect 25872 19246 25924 19252
rect 25780 19236 25832 19242
rect 25780 19178 25832 19184
rect 25320 18692 25372 18698
rect 25320 18634 25372 18640
rect 25332 18426 25360 18634
rect 25320 18420 25372 18426
rect 25320 18362 25372 18368
rect 25792 18222 25820 19178
rect 26056 18284 26108 18290
rect 26056 18226 26108 18232
rect 25320 18216 25372 18222
rect 25320 18158 25372 18164
rect 25504 18216 25556 18222
rect 25504 18158 25556 18164
rect 25780 18216 25832 18222
rect 25780 18158 25832 18164
rect 25136 17740 25188 17746
rect 25136 17682 25188 17688
rect 25228 17740 25280 17746
rect 25228 17682 25280 17688
rect 24860 17604 24912 17610
rect 24860 17546 24912 17552
rect 24768 17536 24820 17542
rect 24768 17478 24820 17484
rect 23664 17332 23716 17338
rect 23664 17274 23716 17280
rect 23480 17060 23532 17066
rect 23480 17002 23532 17008
rect 24584 17060 24636 17066
rect 24584 17002 24636 17008
rect 23388 16720 23440 16726
rect 23388 16662 23440 16668
rect 23112 16516 23164 16522
rect 23112 16458 23164 16464
rect 23124 15910 23152 16458
rect 23400 16046 23428 16662
rect 23492 16658 23520 17002
rect 24216 16992 24268 16998
rect 24216 16934 24268 16940
rect 23480 16652 23532 16658
rect 23480 16594 23532 16600
rect 24228 16590 24256 16934
rect 24216 16584 24268 16590
rect 24216 16526 24268 16532
rect 24492 16516 24544 16522
rect 24492 16458 24544 16464
rect 23480 16176 23532 16182
rect 23480 16118 23532 16124
rect 23388 16040 23440 16046
rect 23388 15982 23440 15988
rect 23112 15904 23164 15910
rect 23112 15846 23164 15852
rect 22652 15564 22704 15570
rect 22652 15506 22704 15512
rect 22652 15428 22704 15434
rect 22652 15370 22704 15376
rect 22664 15162 22692 15370
rect 22652 15156 22704 15162
rect 22652 15098 22704 15104
rect 22008 15020 22060 15026
rect 22008 14962 22060 14968
rect 21640 14476 21692 14482
rect 21640 14418 21692 14424
rect 21548 14408 21600 14414
rect 21548 14350 21600 14356
rect 21560 14074 21588 14350
rect 21548 14068 21600 14074
rect 21548 14010 21600 14016
rect 22020 13938 22048 14962
rect 22928 14952 22980 14958
rect 22928 14894 22980 14900
rect 22940 14482 22968 14894
rect 22192 14476 22244 14482
rect 22192 14418 22244 14424
rect 22928 14476 22980 14482
rect 22928 14418 22980 14424
rect 22008 13932 22060 13938
rect 22008 13874 22060 13880
rect 22020 13818 22048 13874
rect 22020 13790 22140 13818
rect 21456 13184 21508 13190
rect 21456 13126 21508 13132
rect 21468 12170 21496 13126
rect 22112 12850 22140 13790
rect 22100 12844 22152 12850
rect 22100 12786 22152 12792
rect 22204 12322 22232 14418
rect 23400 13734 23428 15982
rect 23492 15706 23520 16118
rect 23480 15700 23532 15706
rect 23480 15642 23532 15648
rect 23492 14074 23520 15642
rect 23848 15632 23900 15638
rect 23848 15574 23900 15580
rect 23572 14408 23624 14414
rect 23572 14350 23624 14356
rect 23480 14068 23532 14074
rect 23480 14010 23532 14016
rect 23584 13870 23612 14350
rect 23572 13864 23624 13870
rect 23572 13806 23624 13812
rect 23860 13802 23888 15574
rect 24032 14952 24084 14958
rect 24032 14894 24084 14900
rect 24044 14618 24072 14894
rect 24032 14612 24084 14618
rect 24032 14554 24084 14560
rect 24044 14006 24072 14554
rect 24032 14000 24084 14006
rect 24032 13942 24084 13948
rect 23848 13796 23900 13802
rect 23848 13738 23900 13744
rect 23388 13728 23440 13734
rect 23388 13670 23440 13676
rect 23400 13394 23428 13670
rect 23112 13388 23164 13394
rect 23112 13330 23164 13336
rect 23388 13388 23440 13394
rect 23388 13330 23440 13336
rect 22836 13184 22888 13190
rect 22836 13126 22888 13132
rect 22928 13184 22980 13190
rect 22928 13126 22980 13132
rect 22848 12986 22876 13126
rect 22836 12980 22888 12986
rect 22836 12922 22888 12928
rect 22940 12918 22968 13126
rect 22928 12912 22980 12918
rect 22928 12854 22980 12860
rect 22836 12844 22888 12850
rect 22836 12786 22888 12792
rect 22376 12640 22428 12646
rect 22376 12582 22428 12588
rect 22112 12306 22232 12322
rect 22100 12300 22232 12306
rect 22152 12294 22232 12300
rect 22100 12242 22152 12248
rect 21456 12164 21508 12170
rect 21456 12106 21508 12112
rect 22204 11830 22232 12294
rect 22388 12170 22416 12582
rect 22376 12164 22428 12170
rect 22376 12106 22428 12112
rect 22192 11824 22244 11830
rect 22192 11766 22244 11772
rect 22284 11688 22336 11694
rect 22284 11630 22336 11636
rect 22296 11354 22324 11630
rect 22284 11348 22336 11354
rect 22284 11290 22336 11296
rect 22848 11150 22876 12786
rect 22940 12442 22968 12854
rect 22928 12436 22980 12442
rect 22928 12378 22980 12384
rect 23124 12306 23152 13330
rect 23664 13184 23716 13190
rect 23664 13126 23716 13132
rect 23676 12986 23704 13126
rect 23664 12980 23716 12986
rect 23664 12922 23716 12928
rect 23860 12782 23888 13738
rect 24044 12850 24072 13942
rect 24032 12844 24084 12850
rect 24032 12786 24084 12792
rect 23848 12776 23900 12782
rect 23848 12718 23900 12724
rect 24400 12640 24452 12646
rect 24400 12582 24452 12588
rect 23112 12300 23164 12306
rect 23112 12242 23164 12248
rect 24412 12238 24440 12582
rect 24400 12232 24452 12238
rect 24400 12174 24452 12180
rect 24032 12164 24084 12170
rect 24032 12106 24084 12112
rect 23296 12096 23348 12102
rect 23296 12038 23348 12044
rect 23756 12096 23808 12102
rect 23756 12038 23808 12044
rect 23020 11824 23072 11830
rect 23020 11766 23072 11772
rect 23032 11354 23060 11766
rect 23020 11348 23072 11354
rect 23020 11290 23072 11296
rect 23308 11218 23336 12038
rect 23768 11694 23796 12038
rect 23756 11688 23808 11694
rect 23756 11630 23808 11636
rect 23848 11552 23900 11558
rect 23848 11494 23900 11500
rect 23296 11212 23348 11218
rect 23296 11154 23348 11160
rect 23860 11150 23888 11494
rect 24044 11354 24072 12106
rect 24308 11552 24360 11558
rect 24308 11494 24360 11500
rect 24032 11348 24084 11354
rect 24032 11290 24084 11296
rect 22836 11144 22888 11150
rect 22836 11086 22888 11092
rect 23848 11144 23900 11150
rect 23848 11086 23900 11092
rect 22560 10464 22612 10470
rect 22560 10406 22612 10412
rect 22572 9994 22600 10406
rect 22560 9988 22612 9994
rect 22560 9930 22612 9936
rect 22848 9654 22876 11086
rect 24320 10742 24348 11494
rect 24308 10736 24360 10742
rect 24308 10678 24360 10684
rect 23112 10464 23164 10470
rect 23112 10406 23164 10412
rect 22836 9648 22888 9654
rect 22836 9590 22888 9596
rect 22836 9512 22888 9518
rect 22836 9454 22888 9460
rect 22848 8838 22876 9454
rect 22284 8832 22336 8838
rect 22284 8774 22336 8780
rect 22836 8832 22888 8838
rect 22836 8774 22888 8780
rect 21456 8356 21508 8362
rect 21456 8298 21508 8304
rect 21364 3188 21416 3194
rect 21364 3130 21416 3136
rect 20588 3012 20668 3040
rect 20536 2994 20588 3000
rect 19720 2650 19748 2994
rect 18696 2644 18748 2650
rect 18696 2586 18748 2592
rect 19708 2644 19760 2650
rect 19708 2586 19760 2592
rect 20548 2514 20576 2994
rect 20536 2508 20588 2514
rect 20536 2450 20588 2456
rect 21468 2446 21496 8298
rect 22008 4480 22060 4486
rect 22008 4422 22060 4428
rect 22020 4214 22048 4422
rect 22008 4208 22060 4214
rect 22008 4150 22060 4156
rect 22008 4072 22060 4078
rect 22008 4014 22060 4020
rect 22020 3602 22048 4014
rect 22008 3596 22060 3602
rect 22008 3538 22060 3544
rect 22192 3596 22244 3602
rect 22192 3538 22244 3544
rect 21916 3460 21968 3466
rect 21916 3402 21968 3408
rect 21928 2650 21956 3402
rect 22008 3392 22060 3398
rect 22008 3334 22060 3340
rect 21916 2644 21968 2650
rect 21916 2586 21968 2592
rect 21456 2440 21508 2446
rect 21456 2382 21508 2388
rect 22020 2378 22048 3334
rect 22204 3126 22232 3538
rect 22192 3120 22244 3126
rect 22192 3062 22244 3068
rect 22296 2530 22324 8774
rect 22376 4684 22428 4690
rect 22376 4626 22428 4632
rect 22652 4684 22704 4690
rect 22652 4626 22704 4632
rect 22388 4570 22416 4626
rect 22388 4542 22600 4570
rect 22572 3670 22600 4542
rect 22560 3664 22612 3670
rect 22560 3606 22612 3612
rect 22572 3126 22600 3606
rect 22560 3120 22612 3126
rect 22560 3062 22612 3068
rect 22664 2990 22692 4626
rect 22928 4480 22980 4486
rect 22928 4422 22980 4428
rect 22940 4078 22968 4422
rect 23124 4282 23152 10406
rect 23664 10056 23716 10062
rect 23664 9998 23716 10004
rect 23676 9654 23704 9998
rect 23664 9648 23716 9654
rect 23664 9590 23716 9596
rect 23848 4616 23900 4622
rect 23848 4558 23900 4564
rect 23296 4548 23348 4554
rect 23296 4490 23348 4496
rect 23112 4276 23164 4282
rect 23112 4218 23164 4224
rect 22928 4072 22980 4078
rect 22928 4014 22980 4020
rect 22940 3534 22968 4014
rect 23020 3936 23072 3942
rect 23020 3878 23072 3884
rect 22928 3528 22980 3534
rect 22928 3470 22980 3476
rect 22652 2984 22704 2990
rect 22652 2926 22704 2932
rect 22112 2514 22324 2530
rect 22100 2508 22336 2514
rect 22152 2502 22284 2508
rect 22100 2450 22152 2456
rect 22284 2450 22336 2456
rect 22940 2378 22968 3470
rect 23032 2922 23060 3878
rect 23124 3738 23152 4218
rect 23308 4010 23336 4490
rect 23388 4140 23440 4146
rect 23388 4082 23440 4088
rect 23296 4004 23348 4010
rect 23296 3946 23348 3952
rect 23400 3738 23428 4082
rect 23112 3732 23164 3738
rect 23112 3674 23164 3680
rect 23388 3732 23440 3738
rect 23388 3674 23440 3680
rect 23124 3602 23152 3674
rect 23112 3596 23164 3602
rect 23112 3538 23164 3544
rect 23860 3534 23888 4558
rect 23848 3528 23900 3534
rect 23848 3470 23900 3476
rect 23020 2916 23072 2922
rect 23020 2858 23072 2864
rect 23032 2446 23060 2858
rect 23480 2508 23532 2514
rect 23480 2450 23532 2456
rect 23020 2440 23072 2446
rect 23020 2382 23072 2388
rect 18052 2372 18104 2378
rect 18052 2314 18104 2320
rect 22008 2372 22060 2378
rect 22008 2314 22060 2320
rect 22928 2372 22980 2378
rect 22928 2314 22980 2320
rect 17960 2304 18012 2310
rect 17960 2246 18012 2252
rect 15212 1414 15332 1442
rect 15212 800 15240 1414
rect 17972 800 18000 2246
rect 18064 1970 18092 2314
rect 20444 2304 20496 2310
rect 20444 2246 20496 2252
rect 20720 2304 20772 2310
rect 20720 2246 20772 2252
rect 20456 2106 20484 2246
rect 20444 2100 20496 2106
rect 20444 2042 20496 2048
rect 18052 1964 18104 1970
rect 18052 1906 18104 1912
rect 20732 800 20760 2246
rect 23492 800 23520 2450
rect 24504 2378 24532 16458
rect 24596 16250 24624 17002
rect 24780 16794 24808 17478
rect 24952 17128 25004 17134
rect 24952 17070 25004 17076
rect 24768 16788 24820 16794
rect 24768 16730 24820 16736
rect 24964 16726 24992 17070
rect 25240 16998 25268 17682
rect 25332 17610 25360 18158
rect 25412 17672 25464 17678
rect 25412 17614 25464 17620
rect 25320 17604 25372 17610
rect 25320 17546 25372 17552
rect 25424 17338 25452 17614
rect 25412 17332 25464 17338
rect 25412 17274 25464 17280
rect 25516 17134 25544 18158
rect 26068 17882 26096 18226
rect 26056 17876 26108 17882
rect 26056 17818 26108 17824
rect 26436 17678 26464 19314
rect 26804 18766 26832 19654
rect 26792 18760 26844 18766
rect 26792 18702 26844 18708
rect 26792 18284 26844 18290
rect 26792 18226 26844 18232
rect 26700 18080 26752 18086
rect 26700 18022 26752 18028
rect 26712 17746 26740 18022
rect 26700 17740 26752 17746
rect 26700 17682 26752 17688
rect 26424 17672 26476 17678
rect 26424 17614 26476 17620
rect 25504 17128 25556 17134
rect 25504 17070 25556 17076
rect 25228 16992 25280 16998
rect 25228 16934 25280 16940
rect 25504 16992 25556 16998
rect 25504 16934 25556 16940
rect 24952 16720 25004 16726
rect 24780 16668 24952 16674
rect 24780 16662 25004 16668
rect 24780 16646 24992 16662
rect 24584 16244 24636 16250
rect 24584 16186 24636 16192
rect 24780 16046 24808 16646
rect 25516 16046 25544 16934
rect 26436 16658 26464 17614
rect 26424 16652 26476 16658
rect 26424 16594 26476 16600
rect 25596 16108 25648 16114
rect 25596 16050 25648 16056
rect 24768 16040 24820 16046
rect 24768 15982 24820 15988
rect 25504 16040 25556 16046
rect 25504 15982 25556 15988
rect 25516 15706 25544 15982
rect 25504 15700 25556 15706
rect 25504 15642 25556 15648
rect 25608 15366 25636 16050
rect 25872 15564 25924 15570
rect 25872 15506 25924 15512
rect 25596 15360 25648 15366
rect 25596 15302 25648 15308
rect 24584 15020 24636 15026
rect 24584 14962 24636 14968
rect 24596 13530 24624 14962
rect 24768 14816 24820 14822
rect 24768 14758 24820 14764
rect 24952 14816 25004 14822
rect 24952 14758 25004 14764
rect 24780 14006 24808 14758
rect 24860 14476 24912 14482
rect 24860 14418 24912 14424
rect 24768 14000 24820 14006
rect 24768 13942 24820 13948
rect 24872 13938 24900 14418
rect 24860 13932 24912 13938
rect 24860 13874 24912 13880
rect 24584 13524 24636 13530
rect 24584 13466 24636 13472
rect 24584 12776 24636 12782
rect 24584 12718 24636 12724
rect 24596 12374 24624 12718
rect 24584 12368 24636 12374
rect 24584 12310 24636 12316
rect 24596 11898 24624 12310
rect 24872 12306 24900 13874
rect 24964 13326 24992 14758
rect 25608 14618 25636 15302
rect 25596 14612 25648 14618
rect 25596 14554 25648 14560
rect 25228 14340 25280 14346
rect 25228 14282 25280 14288
rect 25240 13462 25268 14282
rect 25228 13456 25280 13462
rect 25228 13398 25280 13404
rect 24952 13320 25004 13326
rect 24952 13262 25004 13268
rect 25884 13258 25912 15506
rect 26436 15314 26464 16594
rect 26608 15904 26660 15910
rect 26608 15846 26660 15852
rect 26620 15434 26648 15846
rect 26608 15428 26660 15434
rect 26608 15370 26660 15376
rect 26436 15286 26556 15314
rect 26528 15094 26556 15286
rect 26424 15088 26476 15094
rect 26424 15030 26476 15036
rect 26516 15088 26568 15094
rect 26516 15030 26568 15036
rect 26332 14884 26384 14890
rect 26332 14826 26384 14832
rect 26344 13530 26372 14826
rect 26332 13524 26384 13530
rect 26332 13466 26384 13472
rect 26344 13410 26372 13466
rect 26252 13382 26372 13410
rect 25872 13252 25924 13258
rect 25872 13194 25924 13200
rect 25044 13184 25096 13190
rect 25044 13126 25096 13132
rect 25056 12918 25084 13126
rect 25884 12986 25912 13194
rect 25872 12980 25924 12986
rect 25872 12922 25924 12928
rect 25044 12912 25096 12918
rect 25044 12854 25096 12860
rect 24952 12844 25004 12850
rect 24952 12786 25004 12792
rect 26056 12844 26108 12850
rect 26056 12786 26108 12792
rect 24768 12300 24820 12306
rect 24768 12242 24820 12248
rect 24860 12300 24912 12306
rect 24860 12242 24912 12248
rect 24584 11892 24636 11898
rect 24584 11834 24636 11840
rect 24780 11830 24808 12242
rect 24768 11824 24820 11830
rect 24768 11766 24820 11772
rect 24676 11688 24728 11694
rect 24676 11630 24728 11636
rect 24584 11212 24636 11218
rect 24584 11154 24636 11160
rect 24596 10674 24624 11154
rect 24688 11082 24716 11630
rect 24676 11076 24728 11082
rect 24676 11018 24728 11024
rect 24780 10810 24808 11766
rect 24964 11286 24992 12786
rect 25320 11756 25372 11762
rect 25320 11698 25372 11704
rect 25332 11354 25360 11698
rect 25596 11688 25648 11694
rect 25596 11630 25648 11636
rect 25320 11348 25372 11354
rect 25320 11290 25372 11296
rect 24952 11280 25004 11286
rect 24952 11222 25004 11228
rect 25608 11082 25636 11630
rect 25596 11076 25648 11082
rect 25596 11018 25648 11024
rect 24768 10804 24820 10810
rect 24768 10746 24820 10752
rect 24584 10668 24636 10674
rect 24584 10610 24636 10616
rect 24952 10464 25004 10470
rect 24952 10406 25004 10412
rect 24584 10124 24636 10130
rect 24584 10066 24636 10072
rect 24596 9042 24624 10066
rect 24860 9988 24912 9994
rect 24860 9930 24912 9936
rect 24872 9450 24900 9930
rect 24964 9586 24992 10406
rect 25608 10266 25636 11018
rect 26068 10674 26096 12786
rect 26148 11756 26200 11762
rect 26148 11698 26200 11704
rect 26160 11082 26188 11698
rect 26252 11694 26280 13382
rect 26332 13252 26384 13258
rect 26332 13194 26384 13200
rect 26240 11688 26292 11694
rect 26240 11630 26292 11636
rect 26148 11076 26200 11082
rect 26148 11018 26200 11024
rect 26240 11008 26292 11014
rect 26240 10950 26292 10956
rect 26252 10810 26280 10950
rect 26240 10804 26292 10810
rect 26240 10746 26292 10752
rect 26056 10668 26108 10674
rect 26056 10610 26108 10616
rect 25964 10600 26016 10606
rect 25964 10542 26016 10548
rect 26240 10600 26292 10606
rect 26240 10542 26292 10548
rect 25596 10260 25648 10266
rect 25596 10202 25648 10208
rect 25976 10198 26004 10542
rect 25964 10192 26016 10198
rect 25964 10134 26016 10140
rect 25504 9988 25556 9994
rect 25504 9930 25556 9936
rect 25516 9654 25544 9930
rect 25504 9648 25556 9654
rect 25504 9590 25556 9596
rect 26252 9586 26280 10542
rect 24952 9580 25004 9586
rect 24952 9522 25004 9528
rect 26240 9580 26292 9586
rect 26240 9522 26292 9528
rect 26344 9466 26372 13194
rect 26436 10062 26464 15030
rect 26528 14482 26556 15030
rect 26700 15020 26752 15026
rect 26700 14962 26752 14968
rect 26516 14476 26568 14482
rect 26516 14418 26568 14424
rect 26712 14278 26740 14962
rect 26700 14272 26752 14278
rect 26700 14214 26752 14220
rect 26712 14074 26740 14214
rect 26700 14068 26752 14074
rect 26700 14010 26752 14016
rect 26608 13864 26660 13870
rect 26608 13806 26660 13812
rect 26620 13326 26648 13806
rect 26608 13320 26660 13326
rect 26608 13262 26660 13268
rect 26804 13258 26832 18226
rect 26792 13252 26844 13258
rect 26792 13194 26844 13200
rect 26896 12434 26924 24806
rect 27068 24812 27120 24818
rect 27068 24754 27120 24760
rect 27080 24410 27108 24754
rect 27172 24614 27200 25350
rect 27160 24608 27212 24614
rect 27160 24550 27212 24556
rect 27068 24404 27120 24410
rect 27068 24346 27120 24352
rect 27172 23662 27200 24550
rect 27160 23656 27212 23662
rect 27160 23598 27212 23604
rect 27172 22574 27200 23598
rect 27160 22568 27212 22574
rect 27160 22510 27212 22516
rect 26976 21888 27028 21894
rect 26976 21830 27028 21836
rect 26988 21622 27016 21830
rect 26976 21616 27028 21622
rect 26976 21558 27028 21564
rect 27172 21554 27200 22510
rect 27264 21690 27292 30194
rect 27632 30122 27660 30670
rect 27620 30116 27672 30122
rect 27620 30058 27672 30064
rect 27436 29844 27488 29850
rect 27436 29786 27488 29792
rect 27448 29170 27476 29786
rect 27724 29782 27752 32166
rect 27896 31884 27948 31890
rect 27896 31826 27948 31832
rect 27908 31142 27936 31826
rect 28080 31816 28132 31822
rect 28080 31758 28132 31764
rect 27988 31340 28040 31346
rect 27988 31282 28040 31288
rect 27896 31136 27948 31142
rect 27896 31078 27948 31084
rect 28000 30938 28028 31282
rect 27988 30932 28040 30938
rect 27988 30874 28040 30880
rect 28092 30870 28120 31758
rect 28172 31748 28224 31754
rect 28172 31690 28224 31696
rect 28080 30864 28132 30870
rect 28080 30806 28132 30812
rect 27896 30728 27948 30734
rect 27896 30670 27948 30676
rect 27988 30728 28040 30734
rect 27988 30670 28040 30676
rect 27804 30592 27856 30598
rect 27804 30534 27856 30540
rect 27712 29776 27764 29782
rect 27712 29718 27764 29724
rect 27816 29646 27844 30534
rect 27908 30122 27936 30670
rect 27896 30116 27948 30122
rect 27896 30058 27948 30064
rect 27908 29646 27936 30058
rect 28000 29714 28028 30670
rect 28184 30376 28212 31690
rect 28092 30348 28212 30376
rect 28092 30054 28120 30348
rect 28172 30252 28224 30258
rect 28172 30194 28224 30200
rect 28080 30048 28132 30054
rect 28080 29990 28132 29996
rect 27988 29708 28040 29714
rect 27988 29650 28040 29656
rect 27804 29640 27856 29646
rect 27804 29582 27856 29588
rect 27896 29640 27948 29646
rect 27896 29582 27948 29588
rect 27436 29164 27488 29170
rect 27436 29106 27488 29112
rect 27528 27872 27580 27878
rect 27528 27814 27580 27820
rect 27540 27402 27568 27814
rect 27436 27396 27488 27402
rect 27436 27338 27488 27344
rect 27528 27396 27580 27402
rect 27528 27338 27580 27344
rect 27448 27130 27476 27338
rect 27436 27124 27488 27130
rect 27436 27066 27488 27072
rect 27344 26920 27396 26926
rect 27344 26862 27396 26868
rect 27356 26382 27384 26862
rect 27344 26376 27396 26382
rect 27396 26336 27476 26364
rect 27344 26318 27396 26324
rect 27448 24818 27476 26336
rect 27712 26240 27764 26246
rect 27712 26182 27764 26188
rect 27724 25974 27752 26182
rect 27712 25968 27764 25974
rect 27712 25910 27764 25916
rect 27896 25968 27948 25974
rect 27896 25910 27948 25916
rect 27908 24818 27936 25910
rect 27436 24812 27488 24818
rect 27436 24754 27488 24760
rect 27896 24812 27948 24818
rect 27896 24754 27948 24760
rect 27896 23792 27948 23798
rect 27896 23734 27948 23740
rect 27436 23656 27488 23662
rect 27436 23598 27488 23604
rect 27448 23322 27476 23598
rect 27908 23322 27936 23734
rect 27436 23316 27488 23322
rect 27436 23258 27488 23264
rect 27896 23316 27948 23322
rect 27896 23258 27948 23264
rect 27712 23112 27764 23118
rect 27712 23054 27764 23060
rect 27724 22030 27752 23054
rect 28000 22982 28028 29650
rect 28080 29572 28132 29578
rect 28080 29514 28132 29520
rect 28092 23866 28120 29514
rect 28080 23860 28132 23866
rect 28080 23802 28132 23808
rect 27988 22976 28040 22982
rect 27988 22918 28040 22924
rect 28000 22760 28028 22918
rect 28080 22772 28132 22778
rect 28000 22732 28080 22760
rect 28080 22714 28132 22720
rect 27896 22704 27948 22710
rect 27896 22646 27948 22652
rect 27908 22098 27936 22646
rect 27896 22092 27948 22098
rect 27896 22034 27948 22040
rect 27712 22024 27764 22030
rect 27712 21966 27764 21972
rect 27252 21684 27304 21690
rect 27252 21626 27304 21632
rect 27160 21548 27212 21554
rect 27160 21490 27212 21496
rect 27264 20806 27292 21626
rect 27528 21004 27580 21010
rect 27528 20946 27580 20952
rect 27252 20800 27304 20806
rect 27252 20742 27304 20748
rect 27252 20392 27304 20398
rect 27252 20334 27304 20340
rect 26976 20256 27028 20262
rect 26976 20198 27028 20204
rect 26988 19922 27016 20198
rect 26976 19916 27028 19922
rect 26976 19858 27028 19864
rect 27264 19514 27292 20334
rect 27252 19508 27304 19514
rect 27252 19450 27304 19456
rect 26976 19304 27028 19310
rect 26976 19246 27028 19252
rect 26988 18970 27016 19246
rect 26976 18964 27028 18970
rect 26976 18906 27028 18912
rect 27540 18766 27568 20946
rect 27724 20874 27752 21966
rect 27712 20868 27764 20874
rect 27712 20810 27764 20816
rect 28184 20602 28212 30194
rect 28276 29782 28304 32710
rect 28448 31136 28500 31142
rect 28448 31078 28500 31084
rect 28460 30734 28488 31078
rect 28448 30728 28500 30734
rect 28448 30670 28500 30676
rect 28448 30592 28500 30598
rect 28448 30534 28500 30540
rect 28356 30388 28408 30394
rect 28356 30330 28408 30336
rect 28368 30172 28396 30330
rect 28460 30326 28488 30534
rect 28448 30320 28500 30326
rect 28448 30262 28500 30268
rect 28552 30258 28580 33798
rect 28632 32904 28684 32910
rect 28632 32846 28684 32852
rect 28644 31822 28672 32846
rect 28632 31816 28684 31822
rect 28632 31758 28684 31764
rect 28540 30252 28592 30258
rect 28540 30194 28592 30200
rect 28632 30252 28684 30258
rect 28632 30194 28684 30200
rect 28368 30144 28488 30172
rect 28356 30048 28408 30054
rect 28356 29990 28408 29996
rect 28264 29776 28316 29782
rect 28264 29718 28316 29724
rect 28368 29170 28396 29990
rect 28460 29714 28488 30144
rect 28448 29708 28500 29714
rect 28448 29650 28500 29656
rect 28552 29170 28580 30194
rect 28356 29164 28408 29170
rect 28356 29106 28408 29112
rect 28540 29164 28592 29170
rect 28540 29106 28592 29112
rect 28644 29102 28672 30194
rect 28448 29096 28500 29102
rect 28448 29038 28500 29044
rect 28632 29096 28684 29102
rect 28632 29038 28684 29044
rect 28736 29050 28764 38150
rect 29564 37874 29592 38354
rect 29736 38276 29788 38282
rect 29736 38218 29788 38224
rect 29748 38010 29776 38218
rect 29920 38208 29972 38214
rect 29920 38150 29972 38156
rect 30104 38208 30156 38214
rect 30104 38150 30156 38156
rect 29736 38004 29788 38010
rect 29736 37946 29788 37952
rect 29368 37868 29420 37874
rect 29368 37810 29420 37816
rect 29552 37868 29604 37874
rect 29552 37810 29604 37816
rect 29092 37664 29144 37670
rect 29092 37606 29144 37612
rect 28816 37392 28868 37398
rect 28816 37334 28868 37340
rect 28828 37126 28856 37334
rect 29104 37194 29132 37606
rect 29276 37256 29328 37262
rect 29276 37198 29328 37204
rect 29092 37188 29144 37194
rect 29092 37130 29144 37136
rect 28816 37120 28868 37126
rect 28816 37062 28868 37068
rect 28908 37120 28960 37126
rect 29288 37074 29316 37198
rect 29380 37126 29408 37810
rect 29932 37312 29960 38150
rect 30012 37324 30064 37330
rect 29932 37284 30012 37312
rect 30012 37266 30064 37272
rect 28908 37062 28960 37068
rect 28816 35760 28868 35766
rect 28816 35702 28868 35708
rect 28828 35290 28856 35702
rect 28920 35698 28948 37062
rect 29104 37046 29316 37074
rect 29368 37120 29420 37126
rect 29368 37062 29420 37068
rect 29828 37120 29880 37126
rect 29828 37062 29880 37068
rect 29104 36582 29132 37046
rect 29840 36786 29868 37062
rect 29828 36780 29880 36786
rect 29828 36722 29880 36728
rect 29092 36576 29144 36582
rect 29092 36518 29144 36524
rect 29000 36304 29052 36310
rect 29000 36246 29052 36252
rect 29012 35766 29040 36246
rect 29000 35760 29052 35766
rect 29000 35702 29052 35708
rect 28908 35692 28960 35698
rect 28908 35634 28960 35640
rect 29000 35624 29052 35630
rect 29000 35566 29052 35572
rect 28816 35284 28868 35290
rect 28816 35226 28868 35232
rect 29012 34610 29040 35566
rect 29000 34604 29052 34610
rect 29000 34546 29052 34552
rect 29000 33380 29052 33386
rect 29000 33322 29052 33328
rect 29012 32570 29040 33322
rect 29104 32858 29132 36518
rect 29736 36032 29788 36038
rect 29736 35974 29788 35980
rect 29748 35630 29776 35974
rect 29736 35624 29788 35630
rect 29736 35566 29788 35572
rect 29368 35488 29420 35494
rect 29368 35430 29420 35436
rect 29184 33448 29236 33454
rect 29236 33396 29316 33402
rect 29184 33390 29316 33396
rect 29196 33374 29316 33390
rect 29184 33312 29236 33318
rect 29184 33254 29236 33260
rect 29196 32978 29224 33254
rect 29184 32972 29236 32978
rect 29184 32914 29236 32920
rect 29104 32830 29224 32858
rect 29000 32564 29052 32570
rect 29000 32506 29052 32512
rect 29092 31952 29144 31958
rect 29092 31894 29144 31900
rect 29000 31816 29052 31822
rect 29000 31758 29052 31764
rect 29012 31482 29040 31758
rect 29000 31476 29052 31482
rect 29000 31418 29052 31424
rect 28908 30864 28960 30870
rect 28908 30806 28960 30812
rect 28920 30394 28948 30806
rect 29012 30734 29040 31418
rect 29000 30728 29052 30734
rect 29000 30670 29052 30676
rect 28908 30388 28960 30394
rect 28908 30330 28960 30336
rect 28816 30252 28868 30258
rect 28816 30194 28868 30200
rect 28828 29646 28856 30194
rect 29104 30122 29132 31894
rect 28908 30116 28960 30122
rect 28908 30058 28960 30064
rect 29092 30116 29144 30122
rect 29092 30058 29144 30064
rect 28920 29850 28948 30058
rect 28908 29844 28960 29850
rect 28908 29786 28960 29792
rect 29196 29730 29224 32830
rect 29288 32026 29316 33374
rect 29380 32910 29408 35430
rect 29460 34536 29512 34542
rect 29460 34478 29512 34484
rect 29368 32904 29420 32910
rect 29368 32846 29420 32852
rect 29276 32020 29328 32026
rect 29276 31962 29328 31968
rect 29380 31958 29408 32846
rect 29368 31952 29420 31958
rect 29368 31894 29420 31900
rect 29276 31204 29328 31210
rect 29276 31146 29328 31152
rect 29288 30394 29316 31146
rect 29276 30388 29328 30394
rect 29276 30330 29328 30336
rect 29000 29708 29052 29714
rect 29196 29702 29316 29730
rect 29000 29650 29052 29656
rect 28816 29640 28868 29646
rect 28816 29582 28868 29588
rect 28908 29164 28960 29170
rect 28908 29106 28960 29112
rect 28816 29096 28868 29102
rect 28736 29044 28816 29050
rect 28736 29038 28868 29044
rect 28356 28620 28408 28626
rect 28356 28562 28408 28568
rect 28264 28552 28316 28558
rect 28264 28494 28316 28500
rect 28276 28218 28304 28494
rect 28264 28212 28316 28218
rect 28264 28154 28316 28160
rect 28368 27334 28396 28562
rect 28356 27328 28408 27334
rect 28356 27270 28408 27276
rect 28368 26994 28396 27270
rect 28356 26988 28408 26994
rect 28356 26930 28408 26936
rect 28460 26874 28488 29038
rect 28736 29022 28856 29038
rect 28736 28626 28764 29022
rect 28920 28642 28948 29106
rect 29012 28762 29040 29650
rect 29092 29640 29144 29646
rect 29092 29582 29144 29588
rect 29184 29640 29236 29646
rect 29184 29582 29236 29588
rect 29104 28762 29132 29582
rect 29196 29306 29224 29582
rect 29184 29300 29236 29306
rect 29184 29242 29236 29248
rect 29000 28756 29052 28762
rect 29000 28698 29052 28704
rect 29092 28756 29144 28762
rect 29092 28698 29144 28704
rect 29184 28688 29236 28694
rect 28920 28636 29184 28642
rect 28920 28630 29236 28636
rect 28724 28620 28776 28626
rect 28920 28614 29224 28630
rect 28724 28562 28776 28568
rect 28908 28552 28960 28558
rect 28908 28494 28960 28500
rect 28540 28484 28592 28490
rect 28540 28426 28592 28432
rect 28552 26994 28580 28426
rect 28816 28076 28868 28082
rect 28816 28018 28868 28024
rect 28828 27674 28856 28018
rect 28920 28014 28948 28494
rect 28908 28008 28960 28014
rect 28908 27950 28960 27956
rect 28816 27668 28868 27674
rect 28816 27610 28868 27616
rect 28632 27056 28684 27062
rect 28632 26998 28684 27004
rect 28540 26988 28592 26994
rect 28540 26930 28592 26936
rect 28368 26846 28488 26874
rect 28540 26852 28592 26858
rect 28368 26042 28396 26846
rect 28540 26794 28592 26800
rect 28448 26784 28500 26790
rect 28448 26726 28500 26732
rect 28460 26586 28488 26726
rect 28448 26580 28500 26586
rect 28448 26522 28500 26528
rect 28552 26314 28580 26794
rect 28644 26382 28672 26998
rect 28632 26376 28684 26382
rect 28632 26318 28684 26324
rect 28540 26308 28592 26314
rect 28540 26250 28592 26256
rect 28908 26240 28960 26246
rect 28908 26182 28960 26188
rect 28356 26036 28408 26042
rect 28356 25978 28408 25984
rect 28368 25498 28396 25978
rect 28356 25492 28408 25498
rect 28356 25434 28408 25440
rect 28368 24206 28396 25434
rect 28920 24954 28948 26182
rect 29012 25702 29040 28614
rect 29288 28490 29316 29702
rect 29472 28966 29500 34478
rect 29644 33380 29696 33386
rect 29644 33322 29696 33328
rect 29552 32564 29604 32570
rect 29552 32506 29604 32512
rect 29564 31822 29592 32506
rect 29656 32502 29684 33322
rect 29644 32496 29696 32502
rect 29644 32438 29696 32444
rect 29552 31816 29604 31822
rect 29552 31758 29604 31764
rect 29736 31680 29788 31686
rect 29736 31622 29788 31628
rect 29748 30938 29776 31622
rect 29736 30932 29788 30938
rect 29736 30874 29788 30880
rect 29748 30054 29776 30874
rect 29736 30048 29788 30054
rect 29736 29990 29788 29996
rect 29840 29646 29868 36722
rect 30024 36650 30052 37266
rect 30116 36718 30144 38150
rect 30300 37670 30328 38490
rect 30288 37664 30340 37670
rect 30288 37606 30340 37612
rect 30300 36786 30328 37606
rect 30380 37188 30432 37194
rect 30380 37130 30432 37136
rect 30288 36780 30340 36786
rect 30288 36722 30340 36728
rect 30104 36712 30156 36718
rect 30104 36654 30156 36660
rect 30012 36644 30064 36650
rect 30012 36586 30064 36592
rect 29920 35760 29972 35766
rect 29920 35702 29972 35708
rect 29932 35290 29960 35702
rect 30024 35476 30052 36586
rect 30300 36378 30328 36722
rect 30392 36718 30420 37130
rect 30380 36712 30432 36718
rect 30380 36654 30432 36660
rect 30288 36372 30340 36378
rect 30288 36314 30340 36320
rect 30564 36168 30616 36174
rect 30564 36110 30616 36116
rect 30840 36168 30892 36174
rect 30840 36110 30892 36116
rect 30288 36100 30340 36106
rect 30288 36042 30340 36048
rect 30104 35488 30156 35494
rect 30024 35448 30104 35476
rect 30104 35430 30156 35436
rect 29920 35284 29972 35290
rect 29920 35226 29972 35232
rect 29932 34746 29960 35226
rect 29920 34740 29972 34746
rect 29920 34682 29972 34688
rect 29920 34604 29972 34610
rect 29920 34546 29972 34552
rect 29932 33862 29960 34546
rect 30300 34474 30328 36042
rect 30380 35760 30432 35766
rect 30380 35702 30432 35708
rect 30392 34542 30420 35702
rect 30576 35630 30604 36110
rect 30852 35698 30880 36110
rect 30840 35692 30892 35698
rect 30840 35634 30892 35640
rect 30564 35624 30616 35630
rect 30564 35566 30616 35572
rect 30932 35624 30984 35630
rect 30932 35566 30984 35572
rect 30576 34950 30604 35566
rect 30564 34944 30616 34950
rect 30564 34886 30616 34892
rect 30380 34536 30432 34542
rect 30380 34478 30432 34484
rect 30472 34536 30524 34542
rect 30472 34478 30524 34484
rect 30288 34468 30340 34474
rect 30288 34410 30340 34416
rect 29920 33856 29972 33862
rect 29920 33798 29972 33804
rect 30104 33856 30156 33862
rect 30104 33798 30156 33804
rect 30116 33658 30144 33798
rect 30104 33652 30156 33658
rect 30104 33594 30156 33600
rect 30012 33516 30064 33522
rect 30012 33458 30064 33464
rect 29920 33448 29972 33454
rect 29920 33390 29972 33396
rect 29932 32434 29960 33390
rect 30024 33046 30052 33458
rect 30116 33114 30144 33594
rect 30392 33386 30420 34478
rect 30484 33998 30512 34478
rect 30472 33992 30524 33998
rect 30472 33934 30524 33940
rect 30380 33380 30432 33386
rect 30380 33322 30432 33328
rect 30392 33114 30420 33322
rect 30104 33108 30156 33114
rect 30104 33050 30156 33056
rect 30380 33108 30432 33114
rect 30380 33050 30432 33056
rect 30012 33040 30064 33046
rect 30012 32982 30064 32988
rect 29920 32428 29972 32434
rect 29920 32370 29972 32376
rect 30024 32230 30052 32982
rect 30012 32224 30064 32230
rect 30012 32166 30064 32172
rect 30576 31754 30604 34886
rect 30944 34746 30972 35566
rect 30932 34740 30984 34746
rect 30932 34682 30984 34688
rect 31128 34678 31156 40093
rect 34072 38554 34100 40093
rect 34934 38652 35242 38661
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38587 35242 38596
rect 34060 38548 34112 38554
rect 34060 38490 34112 38496
rect 31392 38344 31444 38350
rect 31392 38286 31444 38292
rect 33508 38344 33560 38350
rect 33508 38286 33560 38292
rect 34704 38344 34756 38350
rect 34704 38286 34756 38292
rect 31300 37324 31352 37330
rect 31300 37266 31352 37272
rect 31208 36372 31260 36378
rect 31208 36314 31260 36320
rect 31220 35766 31248 36314
rect 31312 36242 31340 37266
rect 31404 36922 31432 38286
rect 31484 38208 31536 38214
rect 31484 38150 31536 38156
rect 32404 38208 32456 38214
rect 32404 38150 32456 38156
rect 33048 38208 33100 38214
rect 33048 38150 33100 38156
rect 31496 37942 31524 38150
rect 31484 37936 31536 37942
rect 31484 37878 31536 37884
rect 31760 37800 31812 37806
rect 31760 37742 31812 37748
rect 31772 37330 31800 37742
rect 31760 37324 31812 37330
rect 31760 37266 31812 37272
rect 32416 37262 32444 38150
rect 33060 37942 33088 38150
rect 33416 38004 33468 38010
rect 33416 37946 33468 37952
rect 33048 37936 33100 37942
rect 33048 37878 33100 37884
rect 33428 37262 33456 37946
rect 33520 37262 33548 38286
rect 34716 38010 34744 38286
rect 35594 38108 35902 38117
rect 35594 38106 35600 38108
rect 35656 38106 35680 38108
rect 35736 38106 35760 38108
rect 35816 38106 35840 38108
rect 35896 38106 35902 38108
rect 35656 38054 35658 38106
rect 35838 38054 35840 38106
rect 35594 38052 35600 38054
rect 35656 38052 35680 38054
rect 35736 38052 35760 38054
rect 35816 38052 35840 38054
rect 35896 38052 35902 38054
rect 35594 38043 35902 38052
rect 34704 38004 34756 38010
rect 34704 37946 34756 37952
rect 34520 37868 34572 37874
rect 34520 37810 34572 37816
rect 33784 37800 33836 37806
rect 33784 37742 33836 37748
rect 34060 37800 34112 37806
rect 34060 37742 34112 37748
rect 33796 37466 33824 37742
rect 34072 37670 34100 37742
rect 34060 37664 34112 37670
rect 34060 37606 34112 37612
rect 33784 37460 33836 37466
rect 33784 37402 33836 37408
rect 32404 37256 32456 37262
rect 32404 37198 32456 37204
rect 33416 37256 33468 37262
rect 33416 37198 33468 37204
rect 33508 37256 33560 37262
rect 33508 37198 33560 37204
rect 31392 36916 31444 36922
rect 31392 36858 31444 36864
rect 31300 36236 31352 36242
rect 31300 36178 31352 36184
rect 32312 36236 32364 36242
rect 32312 36178 32364 36184
rect 31668 36032 31720 36038
rect 31668 35974 31720 35980
rect 31208 35760 31260 35766
rect 31208 35702 31260 35708
rect 31116 34672 31168 34678
rect 31116 34614 31168 34620
rect 31220 34610 31248 35702
rect 31484 35488 31536 35494
rect 31484 35430 31536 35436
rect 31496 34610 31524 35430
rect 31680 34610 31708 35974
rect 32324 35698 32352 36178
rect 33520 36174 33548 37198
rect 34072 36854 34100 37606
rect 34060 36848 34112 36854
rect 34060 36790 34112 36796
rect 33600 36780 33652 36786
rect 33600 36722 33652 36728
rect 33508 36168 33560 36174
rect 33508 36110 33560 36116
rect 33048 36100 33100 36106
rect 33048 36042 33100 36048
rect 32312 35692 32364 35698
rect 32312 35634 32364 35640
rect 32324 35154 32352 35634
rect 33060 35290 33088 36042
rect 33048 35284 33100 35290
rect 33048 35226 33100 35232
rect 32312 35148 32364 35154
rect 32312 35090 32364 35096
rect 33520 35086 33548 36110
rect 33508 35080 33560 35086
rect 33508 35022 33560 35028
rect 32680 35012 32732 35018
rect 32680 34954 32732 34960
rect 32692 34746 32720 34954
rect 33140 34944 33192 34950
rect 33140 34886 33192 34892
rect 32680 34740 32732 34746
rect 32680 34682 32732 34688
rect 31208 34604 31260 34610
rect 31208 34546 31260 34552
rect 31484 34604 31536 34610
rect 31484 34546 31536 34552
rect 31668 34604 31720 34610
rect 31668 34546 31720 34552
rect 33152 34202 33180 34886
rect 33140 34196 33192 34202
rect 33140 34138 33192 34144
rect 33520 33998 33548 35022
rect 33612 34474 33640 36722
rect 33692 36032 33744 36038
rect 33692 35974 33744 35980
rect 33704 35698 33732 35974
rect 33692 35692 33744 35698
rect 33692 35634 33744 35640
rect 33600 34468 33652 34474
rect 33600 34410 33652 34416
rect 32772 33992 32824 33998
rect 32772 33934 32824 33940
rect 33508 33992 33560 33998
rect 33508 33934 33560 33940
rect 32404 33924 32456 33930
rect 32404 33866 32456 33872
rect 32416 33658 32444 33866
rect 32404 33652 32456 33658
rect 32404 33594 32456 33600
rect 31392 33516 31444 33522
rect 31392 33458 31444 33464
rect 31404 33046 31432 33458
rect 31300 33040 31352 33046
rect 31300 32982 31352 32988
rect 31392 33040 31444 33046
rect 31392 32982 31444 32988
rect 30932 32564 30984 32570
rect 30932 32506 30984 32512
rect 30840 32224 30892 32230
rect 30840 32166 30892 32172
rect 30748 31884 30800 31890
rect 30748 31826 30800 31832
rect 30656 31816 30708 31822
rect 30656 31758 30708 31764
rect 30484 31726 30604 31754
rect 29920 31680 29972 31686
rect 29920 31622 29972 31628
rect 29932 30802 29960 31622
rect 29920 30796 29972 30802
rect 29920 30738 29972 30744
rect 29920 29776 29972 29782
rect 29920 29718 29972 29724
rect 29552 29640 29604 29646
rect 29552 29582 29604 29588
rect 29828 29640 29880 29646
rect 29828 29582 29880 29588
rect 29564 29306 29592 29582
rect 29736 29504 29788 29510
rect 29736 29446 29788 29452
rect 29552 29300 29604 29306
rect 29552 29242 29604 29248
rect 29644 29300 29696 29306
rect 29644 29242 29696 29248
rect 29460 28960 29512 28966
rect 29460 28902 29512 28908
rect 29472 28490 29500 28902
rect 29656 28626 29684 29242
rect 29644 28620 29696 28626
rect 29644 28562 29696 28568
rect 29276 28484 29328 28490
rect 29276 28426 29328 28432
rect 29460 28484 29512 28490
rect 29460 28426 29512 28432
rect 29184 27872 29236 27878
rect 29184 27814 29236 27820
rect 29196 27130 29224 27814
rect 29184 27124 29236 27130
rect 29184 27066 29236 27072
rect 29276 26784 29328 26790
rect 29276 26726 29328 26732
rect 29000 25696 29052 25702
rect 29000 25638 29052 25644
rect 29288 25226 29316 26726
rect 29748 25906 29776 29446
rect 29840 29170 29868 29582
rect 29828 29164 29880 29170
rect 29828 29106 29880 29112
rect 29828 28552 29880 28558
rect 29828 28494 29880 28500
rect 29840 27878 29868 28494
rect 29932 28422 29960 29718
rect 30012 29572 30064 29578
rect 30012 29514 30064 29520
rect 30024 29238 30052 29514
rect 30012 29232 30064 29238
rect 30012 29174 30064 29180
rect 30380 29096 30432 29102
rect 30380 29038 30432 29044
rect 29920 28416 29972 28422
rect 29920 28358 29972 28364
rect 29932 28218 29960 28358
rect 29920 28212 29972 28218
rect 29920 28154 29972 28160
rect 29828 27872 29880 27878
rect 29828 27814 29880 27820
rect 29736 25900 29788 25906
rect 29736 25842 29788 25848
rect 29368 25696 29420 25702
rect 29368 25638 29420 25644
rect 29380 25294 29408 25638
rect 29748 25498 29776 25842
rect 30392 25786 30420 29038
rect 30484 27946 30512 31726
rect 30564 30932 30616 30938
rect 30564 30874 30616 30880
rect 30576 30190 30604 30874
rect 30564 30184 30616 30190
rect 30564 30126 30616 30132
rect 30668 29510 30696 31758
rect 30760 31142 30788 31826
rect 30852 31210 30880 32166
rect 30944 32026 30972 32506
rect 31312 32434 31340 32982
rect 31116 32428 31168 32434
rect 31116 32370 31168 32376
rect 31300 32428 31352 32434
rect 31300 32370 31352 32376
rect 30932 32020 30984 32026
rect 30932 31962 30984 31968
rect 30944 31822 30972 31962
rect 30932 31816 30984 31822
rect 30932 31758 30984 31764
rect 30840 31204 30892 31210
rect 30840 31146 30892 31152
rect 30944 31142 30972 31758
rect 31128 31414 31156 32370
rect 31312 32298 31340 32370
rect 31300 32292 31352 32298
rect 31300 32234 31352 32240
rect 31312 31414 31340 32234
rect 31404 32212 31432 32982
rect 32784 32910 32812 33934
rect 33048 33856 33100 33862
rect 33048 33798 33100 33804
rect 33060 33658 33088 33798
rect 33048 33652 33100 33658
rect 33048 33594 33100 33600
rect 33520 33522 33548 33934
rect 33508 33516 33560 33522
rect 33508 33458 33560 33464
rect 33508 32972 33560 32978
rect 33508 32914 33560 32920
rect 32772 32904 32824 32910
rect 32772 32846 32824 32852
rect 32036 32836 32088 32842
rect 32036 32778 32088 32784
rect 32048 32502 32076 32778
rect 32036 32496 32088 32502
rect 32036 32438 32088 32444
rect 32404 32292 32456 32298
rect 32404 32234 32456 32240
rect 31484 32224 31536 32230
rect 31404 32184 31484 32212
rect 31484 32166 31536 32172
rect 31576 31748 31628 31754
rect 31576 31690 31628 31696
rect 31116 31408 31168 31414
rect 31116 31350 31168 31356
rect 31300 31408 31352 31414
rect 31300 31350 31352 31356
rect 31484 31408 31536 31414
rect 31484 31350 31536 31356
rect 30748 31136 30800 31142
rect 30748 31078 30800 31084
rect 30932 31136 30984 31142
rect 30932 31078 30984 31084
rect 30760 30802 30788 31078
rect 30840 30864 30892 30870
rect 30944 30818 30972 31078
rect 31128 30954 31156 31350
rect 31128 30938 31248 30954
rect 31128 30932 31260 30938
rect 31128 30926 31208 30932
rect 31208 30874 31260 30880
rect 30892 30812 30972 30818
rect 30840 30806 30972 30812
rect 30748 30796 30800 30802
rect 30852 30790 30972 30806
rect 30748 30738 30800 30744
rect 30944 30258 30972 30790
rect 31496 30258 31524 31350
rect 30932 30252 30984 30258
rect 30932 30194 30984 30200
rect 31484 30252 31536 30258
rect 31484 30194 31536 30200
rect 31588 30190 31616 31690
rect 32416 31686 32444 32234
rect 32784 31890 32812 32846
rect 33048 32836 33100 32842
rect 33048 32778 33100 32784
rect 33140 32836 33192 32842
rect 33140 32778 33192 32784
rect 33060 32570 33088 32778
rect 33048 32564 33100 32570
rect 33048 32506 33100 32512
rect 32772 31884 32824 31890
rect 32772 31826 32824 31832
rect 32404 31680 32456 31686
rect 32404 31622 32456 31628
rect 31668 31408 31720 31414
rect 31668 31350 31720 31356
rect 31576 30184 31628 30190
rect 31576 30126 31628 30132
rect 30748 29572 30800 29578
rect 30748 29514 30800 29520
rect 30656 29504 30708 29510
rect 30656 29446 30708 29452
rect 30668 28098 30696 29446
rect 30760 28218 30788 29514
rect 31116 29504 31168 29510
rect 31116 29446 31168 29452
rect 31024 28416 31076 28422
rect 31024 28358 31076 28364
rect 31128 28370 31156 29446
rect 31680 29306 31708 31350
rect 32416 30802 32444 31622
rect 32404 30796 32456 30802
rect 32404 30738 32456 30744
rect 32128 30252 32180 30258
rect 32128 30194 32180 30200
rect 33048 30252 33100 30258
rect 33048 30194 33100 30200
rect 32036 29640 32088 29646
rect 32036 29582 32088 29588
rect 31300 29300 31352 29306
rect 31300 29242 31352 29248
rect 31668 29300 31720 29306
rect 31668 29242 31720 29248
rect 31312 28762 31340 29242
rect 32048 29238 32076 29582
rect 32036 29232 32088 29238
rect 32036 29174 32088 29180
rect 31760 29164 31812 29170
rect 31760 29106 31812 29112
rect 31300 28756 31352 28762
rect 31300 28698 31352 28704
rect 31208 28416 31260 28422
rect 31128 28364 31208 28370
rect 31128 28358 31260 28364
rect 30748 28212 30800 28218
rect 30748 28154 30800 28160
rect 30576 28070 30696 28098
rect 30576 28014 30604 28070
rect 30564 28008 30616 28014
rect 30564 27950 30616 27956
rect 30472 27940 30524 27946
rect 30472 27882 30524 27888
rect 31036 27470 31064 28358
rect 31128 28342 31248 28358
rect 31128 28082 31156 28342
rect 31116 28076 31168 28082
rect 31116 28018 31168 28024
rect 31576 28076 31628 28082
rect 31576 28018 31628 28024
rect 31392 28008 31444 28014
rect 31392 27950 31444 27956
rect 31404 27470 31432 27950
rect 31024 27464 31076 27470
rect 31024 27406 31076 27412
rect 31392 27464 31444 27470
rect 31392 27406 31444 27412
rect 31588 27402 31616 28018
rect 31772 27606 31800 29106
rect 31944 28552 31996 28558
rect 31944 28494 31996 28500
rect 31956 28014 31984 28494
rect 31944 28008 31996 28014
rect 31944 27950 31996 27956
rect 31760 27600 31812 27606
rect 31760 27542 31812 27548
rect 31576 27396 31628 27402
rect 31576 27338 31628 27344
rect 30748 27328 30800 27334
rect 30748 27270 30800 27276
rect 30840 27328 30892 27334
rect 30840 27270 30892 27276
rect 30760 27130 30788 27270
rect 30748 27124 30800 27130
rect 30748 27066 30800 27072
rect 30472 26988 30524 26994
rect 30472 26930 30524 26936
rect 30484 26586 30512 26930
rect 30564 26920 30616 26926
rect 30564 26862 30616 26868
rect 30472 26580 30524 26586
rect 30472 26522 30524 26528
rect 30472 25900 30524 25906
rect 30472 25842 30524 25848
rect 30300 25758 30420 25786
rect 29736 25492 29788 25498
rect 29736 25434 29788 25440
rect 29368 25288 29420 25294
rect 29368 25230 29420 25236
rect 29736 25288 29788 25294
rect 29736 25230 29788 25236
rect 29276 25220 29328 25226
rect 29276 25162 29328 25168
rect 28908 24948 28960 24954
rect 28908 24890 28960 24896
rect 29092 24880 29144 24886
rect 29092 24822 29144 24828
rect 29000 24608 29052 24614
rect 29000 24550 29052 24556
rect 28356 24200 28408 24206
rect 28356 24142 28408 24148
rect 28448 23044 28500 23050
rect 28448 22986 28500 22992
rect 28460 22166 28488 22986
rect 28632 22976 28684 22982
rect 28632 22918 28684 22924
rect 28448 22160 28500 22166
rect 28448 22102 28500 22108
rect 28460 20942 28488 22102
rect 28644 21350 28672 22918
rect 28724 22092 28776 22098
rect 28724 22034 28776 22040
rect 28632 21344 28684 21350
rect 28632 21286 28684 21292
rect 28736 21146 28764 22034
rect 28724 21140 28776 21146
rect 28724 21082 28776 21088
rect 29012 20942 29040 24550
rect 29104 23322 29132 24822
rect 29748 24818 29776 25230
rect 30300 24954 30328 25758
rect 30380 25696 30432 25702
rect 30380 25638 30432 25644
rect 30392 25294 30420 25638
rect 30380 25288 30432 25294
rect 30380 25230 30432 25236
rect 30380 25152 30432 25158
rect 30380 25094 30432 25100
rect 30288 24948 30340 24954
rect 30288 24890 30340 24896
rect 29736 24812 29788 24818
rect 29736 24754 29788 24760
rect 30012 24812 30064 24818
rect 30012 24754 30064 24760
rect 29460 24744 29512 24750
rect 29920 24744 29972 24750
rect 29460 24686 29512 24692
rect 29840 24692 29920 24698
rect 29840 24686 29972 24692
rect 29092 23316 29144 23322
rect 29092 23258 29144 23264
rect 29368 22024 29420 22030
rect 29368 21966 29420 21972
rect 29184 21888 29236 21894
rect 29184 21830 29236 21836
rect 28448 20936 28500 20942
rect 28448 20878 28500 20884
rect 29000 20936 29052 20942
rect 29000 20878 29052 20884
rect 28724 20868 28776 20874
rect 28724 20810 28776 20816
rect 28172 20596 28224 20602
rect 28172 20538 28224 20544
rect 28184 20058 28212 20538
rect 28736 20466 28764 20810
rect 29196 20602 29224 21830
rect 29380 21418 29408 21966
rect 29368 21412 29420 21418
rect 29368 21354 29420 21360
rect 29184 20596 29236 20602
rect 29184 20538 29236 20544
rect 28724 20460 28776 20466
rect 28724 20402 28776 20408
rect 28264 20256 28316 20262
rect 28264 20198 28316 20204
rect 28172 20052 28224 20058
rect 28172 19994 28224 20000
rect 28276 19786 28304 20198
rect 28264 19780 28316 19786
rect 28264 19722 28316 19728
rect 28736 19378 28764 20402
rect 29000 19508 29052 19514
rect 29000 19450 29052 19456
rect 28724 19372 28776 19378
rect 28724 19314 28776 19320
rect 28448 19168 28500 19174
rect 28448 19110 28500 19116
rect 27528 18760 27580 18766
rect 27528 18702 27580 18708
rect 27540 18358 27568 18702
rect 28356 18692 28408 18698
rect 28460 18680 28488 19110
rect 28408 18652 28488 18680
rect 28356 18634 28408 18640
rect 27528 18352 27580 18358
rect 27528 18294 27580 18300
rect 26976 18216 27028 18222
rect 26976 18158 27028 18164
rect 28080 18216 28132 18222
rect 28080 18158 28132 18164
rect 26988 13938 27016 18158
rect 27804 17672 27856 17678
rect 27804 17614 27856 17620
rect 27252 17196 27304 17202
rect 27252 17138 27304 17144
rect 27160 17128 27212 17134
rect 27160 17070 27212 17076
rect 27068 16992 27120 16998
rect 27068 16934 27120 16940
rect 27080 16522 27108 16934
rect 27172 16658 27200 17070
rect 27264 16794 27292 17138
rect 27252 16788 27304 16794
rect 27252 16730 27304 16736
rect 27620 16788 27672 16794
rect 27620 16730 27672 16736
rect 27160 16652 27212 16658
rect 27160 16594 27212 16600
rect 27068 16516 27120 16522
rect 27068 16458 27120 16464
rect 27172 16114 27200 16594
rect 27160 16108 27212 16114
rect 27160 16050 27212 16056
rect 27068 15428 27120 15434
rect 27068 15370 27120 15376
rect 27080 15162 27108 15370
rect 27068 15156 27120 15162
rect 27068 15098 27120 15104
rect 27172 14074 27200 16050
rect 27632 15502 27660 16730
rect 27816 16590 27844 17614
rect 28092 17134 28120 18158
rect 28172 17536 28224 17542
rect 28172 17478 28224 17484
rect 28080 17128 28132 17134
rect 28080 17070 28132 17076
rect 27804 16584 27856 16590
rect 27804 16526 27856 16532
rect 27712 16108 27764 16114
rect 27712 16050 27764 16056
rect 27344 15496 27396 15502
rect 27344 15438 27396 15444
rect 27620 15496 27672 15502
rect 27620 15438 27672 15444
rect 27356 15094 27384 15438
rect 27344 15088 27396 15094
rect 27344 15030 27396 15036
rect 27252 14340 27304 14346
rect 27252 14282 27304 14288
rect 27160 14068 27212 14074
rect 27160 14010 27212 14016
rect 26976 13932 27028 13938
rect 26976 13874 27028 13880
rect 27172 12850 27200 14010
rect 27264 12986 27292 14282
rect 27356 13394 27384 15030
rect 27724 14618 27752 16050
rect 27712 14612 27764 14618
rect 27712 14554 27764 14560
rect 27436 13864 27488 13870
rect 27436 13806 27488 13812
rect 27620 13864 27672 13870
rect 27620 13806 27672 13812
rect 27344 13388 27396 13394
rect 27344 13330 27396 13336
rect 27252 12980 27304 12986
rect 27252 12922 27304 12928
rect 27448 12850 27476 13806
rect 27528 13524 27580 13530
rect 27528 13466 27580 13472
rect 27160 12844 27212 12850
rect 27160 12786 27212 12792
rect 27436 12844 27488 12850
rect 27436 12786 27488 12792
rect 26896 12406 27016 12434
rect 26608 11824 26660 11830
rect 26608 11766 26660 11772
rect 26620 11218 26648 11766
rect 26608 11212 26660 11218
rect 26608 11154 26660 11160
rect 26988 10742 27016 12406
rect 27344 12164 27396 12170
rect 27344 12106 27396 12112
rect 27356 11898 27384 12106
rect 27344 11892 27396 11898
rect 27344 11834 27396 11840
rect 27540 11830 27568 13466
rect 27528 11824 27580 11830
rect 27528 11766 27580 11772
rect 27632 11762 27660 13806
rect 28092 12306 28120 17070
rect 28184 16658 28212 17478
rect 28172 16652 28224 16658
rect 28172 16594 28224 16600
rect 28264 14884 28316 14890
rect 28264 14826 28316 14832
rect 28276 14482 28304 14826
rect 28264 14476 28316 14482
rect 28264 14418 28316 14424
rect 28264 14340 28316 14346
rect 28264 14282 28316 14288
rect 28276 13870 28304 14282
rect 28264 13864 28316 13870
rect 28264 13806 28316 13812
rect 28276 12986 28304 13806
rect 28368 13734 28396 18634
rect 28540 18284 28592 18290
rect 28540 18226 28592 18232
rect 28632 18284 28684 18290
rect 28632 18226 28684 18232
rect 28552 17338 28580 18226
rect 28644 17882 28672 18226
rect 28632 17876 28684 17882
rect 28632 17818 28684 17824
rect 28540 17332 28592 17338
rect 28540 17274 28592 17280
rect 28736 16726 28764 19314
rect 29012 18766 29040 19450
rect 29000 18760 29052 18766
rect 29000 18702 29052 18708
rect 29184 18760 29236 18766
rect 29184 18702 29236 18708
rect 28816 18624 28868 18630
rect 28816 18566 28868 18572
rect 28828 18358 28856 18566
rect 28816 18352 28868 18358
rect 28816 18294 28868 18300
rect 28908 17672 28960 17678
rect 29012 17660 29040 18702
rect 29092 18284 29144 18290
rect 29092 18226 29144 18232
rect 28960 17632 29040 17660
rect 28908 17614 28960 17620
rect 29104 17490 29132 18226
rect 29196 17678 29224 18702
rect 29472 18426 29500 24686
rect 29840 24670 29960 24686
rect 29840 24614 29868 24670
rect 30024 24614 30052 24754
rect 30392 24614 30420 25094
rect 30484 24682 30512 25842
rect 30576 25362 30604 26862
rect 30852 26858 30880 27270
rect 31392 27056 31444 27062
rect 31392 26998 31444 27004
rect 30840 26852 30892 26858
rect 30840 26794 30892 26800
rect 30656 26512 30708 26518
rect 30656 26454 30708 26460
rect 30668 25906 30696 26454
rect 31208 26308 31260 26314
rect 31208 26250 31260 26256
rect 30656 25900 30708 25906
rect 30656 25842 30708 25848
rect 31116 25900 31168 25906
rect 31116 25842 31168 25848
rect 31128 25498 31156 25842
rect 31116 25492 31168 25498
rect 31116 25434 31168 25440
rect 30564 25356 30616 25362
rect 30564 25298 30616 25304
rect 30656 25356 30708 25362
rect 30656 25298 30708 25304
rect 30576 24954 30604 25298
rect 30564 24948 30616 24954
rect 30564 24890 30616 24896
rect 30668 24750 30696 25298
rect 30748 24880 30800 24886
rect 30748 24822 30800 24828
rect 30656 24744 30708 24750
rect 30656 24686 30708 24692
rect 30472 24676 30524 24682
rect 30472 24618 30524 24624
rect 29828 24608 29880 24614
rect 29828 24550 29880 24556
rect 30012 24608 30064 24614
rect 30012 24550 30064 24556
rect 30380 24608 30432 24614
rect 30380 24550 30432 24556
rect 29736 23112 29788 23118
rect 29736 23054 29788 23060
rect 29748 22438 29776 23054
rect 29828 22976 29880 22982
rect 29828 22918 29880 22924
rect 29736 22432 29788 22438
rect 29736 22374 29788 22380
rect 29552 22024 29604 22030
rect 29552 21966 29604 21972
rect 29564 21690 29592 21966
rect 29552 21684 29604 21690
rect 29552 21626 29604 21632
rect 29748 21622 29776 22374
rect 29840 22030 29868 22918
rect 30024 22094 30052 24550
rect 30392 24256 30420 24550
rect 30484 24410 30604 24426
rect 30472 24404 30604 24410
rect 30524 24398 30604 24404
rect 30472 24346 30524 24352
rect 30472 24268 30524 24274
rect 30392 24228 30472 24256
rect 30392 23746 30420 24228
rect 30472 24210 30524 24216
rect 30116 23718 30420 23746
rect 30472 23792 30524 23798
rect 30472 23734 30524 23740
rect 30116 23662 30144 23718
rect 30104 23656 30156 23662
rect 30104 23598 30156 23604
rect 30484 23322 30512 23734
rect 30472 23316 30524 23322
rect 30472 23258 30524 23264
rect 30576 23118 30604 24398
rect 30564 23112 30616 23118
rect 30564 23054 30616 23060
rect 30576 22982 30604 23054
rect 30656 23044 30708 23050
rect 30656 22986 30708 22992
rect 30564 22976 30616 22982
rect 30564 22918 30616 22924
rect 30668 22710 30696 22986
rect 30656 22704 30708 22710
rect 30656 22646 30708 22652
rect 30760 22642 30788 24822
rect 31220 24818 31248 26250
rect 31300 26240 31352 26246
rect 31300 26182 31352 26188
rect 31312 25906 31340 26182
rect 31300 25900 31352 25906
rect 31300 25842 31352 25848
rect 31404 25294 31432 26998
rect 31588 25974 31616 27338
rect 31668 26784 31720 26790
rect 31668 26726 31720 26732
rect 31680 26450 31708 26726
rect 31668 26444 31720 26450
rect 31668 26386 31720 26392
rect 31956 26382 31984 27950
rect 32048 27878 32076 29174
rect 32036 27872 32088 27878
rect 32036 27814 32088 27820
rect 31944 26376 31996 26382
rect 31944 26318 31996 26324
rect 31576 25968 31628 25974
rect 31576 25910 31628 25916
rect 31760 25832 31812 25838
rect 31760 25774 31812 25780
rect 31772 25498 31800 25774
rect 31484 25492 31536 25498
rect 31484 25434 31536 25440
rect 31760 25492 31812 25498
rect 31760 25434 31812 25440
rect 31392 25288 31444 25294
rect 31392 25230 31444 25236
rect 31496 24886 31524 25434
rect 31484 24880 31536 24886
rect 31484 24822 31536 24828
rect 31208 24812 31260 24818
rect 31208 24754 31260 24760
rect 31392 24676 31444 24682
rect 31392 24618 31444 24624
rect 31116 22976 31168 22982
rect 31116 22918 31168 22924
rect 30748 22636 30800 22642
rect 30748 22578 30800 22584
rect 30380 22500 30432 22506
rect 30380 22442 30432 22448
rect 30024 22066 30144 22094
rect 29828 22024 29880 22030
rect 29828 21966 29880 21972
rect 29736 21616 29788 21622
rect 29736 21558 29788 21564
rect 29736 20936 29788 20942
rect 29736 20878 29788 20884
rect 29748 20398 29776 20878
rect 29736 20392 29788 20398
rect 29736 20334 29788 20340
rect 29748 19718 29776 20334
rect 29736 19712 29788 19718
rect 29736 19654 29788 19660
rect 29460 18420 29512 18426
rect 29460 18362 29512 18368
rect 29460 18080 29512 18086
rect 29460 18022 29512 18028
rect 29184 17672 29236 17678
rect 29184 17614 29236 17620
rect 29012 17462 29132 17490
rect 29012 17202 29040 17462
rect 29000 17196 29052 17202
rect 29000 17138 29052 17144
rect 29012 16726 29040 17138
rect 29184 16788 29236 16794
rect 29184 16730 29236 16736
rect 28724 16720 28776 16726
rect 28724 16662 28776 16668
rect 29000 16720 29052 16726
rect 29000 16662 29052 16668
rect 28632 16516 28684 16522
rect 28632 16458 28684 16464
rect 28644 16182 28672 16458
rect 28724 16448 28776 16454
rect 28724 16390 28776 16396
rect 28632 16176 28684 16182
rect 28632 16118 28684 16124
rect 28448 16108 28500 16114
rect 28448 16050 28500 16056
rect 28460 15706 28488 16050
rect 28632 16040 28684 16046
rect 28632 15982 28684 15988
rect 28540 15972 28592 15978
rect 28540 15914 28592 15920
rect 28448 15700 28500 15706
rect 28448 15642 28500 15648
rect 28448 15496 28500 15502
rect 28448 15438 28500 15444
rect 28460 14618 28488 15438
rect 28552 15026 28580 15914
rect 28540 15020 28592 15026
rect 28540 14962 28592 14968
rect 28644 14618 28672 15982
rect 28736 15978 28764 16390
rect 28816 16244 28868 16250
rect 28816 16186 28868 16192
rect 28724 15972 28776 15978
rect 28724 15914 28776 15920
rect 28736 15570 28764 15914
rect 28724 15564 28776 15570
rect 28724 15506 28776 15512
rect 28448 14612 28500 14618
rect 28448 14554 28500 14560
rect 28632 14612 28684 14618
rect 28632 14554 28684 14560
rect 28724 14544 28776 14550
rect 28724 14486 28776 14492
rect 28736 13938 28764 14486
rect 28828 14414 28856 16186
rect 29000 15904 29052 15910
rect 29000 15846 29052 15852
rect 28908 15564 28960 15570
rect 28908 15506 28960 15512
rect 28920 15026 28948 15506
rect 28908 15020 28960 15026
rect 28908 14962 28960 14968
rect 28816 14408 28868 14414
rect 28816 14350 28868 14356
rect 28724 13932 28776 13938
rect 28724 13874 28776 13880
rect 28356 13728 28408 13734
rect 28356 13670 28408 13676
rect 28828 13530 28856 14350
rect 29012 13938 29040 15846
rect 29092 14272 29144 14278
rect 29092 14214 29144 14220
rect 29104 13938 29132 14214
rect 29000 13932 29052 13938
rect 29000 13874 29052 13880
rect 29092 13932 29144 13938
rect 29092 13874 29144 13880
rect 29196 13802 29224 16730
rect 29472 16114 29500 18022
rect 29920 17672 29972 17678
rect 29920 17614 29972 17620
rect 29932 17338 29960 17614
rect 29920 17332 29972 17338
rect 29920 17274 29972 17280
rect 29736 16584 29788 16590
rect 29736 16526 29788 16532
rect 30012 16584 30064 16590
rect 30012 16526 30064 16532
rect 29460 16108 29512 16114
rect 29460 16050 29512 16056
rect 29552 16108 29604 16114
rect 29552 16050 29604 16056
rect 29460 15496 29512 15502
rect 29460 15438 29512 15444
rect 29472 15026 29500 15438
rect 29564 15162 29592 16050
rect 29748 15706 29776 16526
rect 30024 16250 30052 16526
rect 30116 16454 30144 22066
rect 30288 22092 30340 22098
rect 30288 22034 30340 22040
rect 30300 21690 30328 22034
rect 30392 22030 30420 22442
rect 30760 22094 30788 22578
rect 30576 22066 30788 22094
rect 30380 22024 30432 22030
rect 30380 21966 30432 21972
rect 30288 21684 30340 21690
rect 30288 21626 30340 21632
rect 30392 21622 30420 21966
rect 30380 21616 30432 21622
rect 30380 21558 30432 21564
rect 30576 21554 30604 22066
rect 30564 21548 30616 21554
rect 30564 21490 30616 21496
rect 30472 21480 30524 21486
rect 30300 21440 30472 21468
rect 30300 21350 30328 21440
rect 30472 21422 30524 21428
rect 30288 21344 30340 21350
rect 30288 21286 30340 21292
rect 30380 21344 30432 21350
rect 30380 21286 30432 21292
rect 30392 20466 30420 21286
rect 30472 20868 30524 20874
rect 30472 20810 30524 20816
rect 30484 20602 30512 20810
rect 30576 20806 30604 21490
rect 30840 21344 30892 21350
rect 30840 21286 30892 21292
rect 30564 20800 30616 20806
rect 30564 20742 30616 20748
rect 30472 20596 30524 20602
rect 30472 20538 30524 20544
rect 30380 20460 30432 20466
rect 30380 20402 30432 20408
rect 30576 20330 30604 20742
rect 30852 20466 30880 21286
rect 30840 20460 30892 20466
rect 30840 20402 30892 20408
rect 30564 20324 30616 20330
rect 30564 20266 30616 20272
rect 30840 19780 30892 19786
rect 30840 19722 30892 19728
rect 30852 19514 30880 19722
rect 30840 19508 30892 19514
rect 30840 19450 30892 19456
rect 30564 19372 30616 19378
rect 30564 19314 30616 19320
rect 30288 18624 30340 18630
rect 30288 18566 30340 18572
rect 30300 18358 30328 18566
rect 30288 18352 30340 18358
rect 30288 18294 30340 18300
rect 30380 18216 30432 18222
rect 30380 18158 30432 18164
rect 30392 17746 30420 18158
rect 30380 17740 30432 17746
rect 30380 17682 30432 17688
rect 30288 17536 30340 17542
rect 30288 17478 30340 17484
rect 30392 17490 30420 17682
rect 30300 17270 30328 17478
rect 30392 17462 30512 17490
rect 30380 17332 30432 17338
rect 30380 17274 30432 17280
rect 30288 17264 30340 17270
rect 30288 17206 30340 17212
rect 30104 16448 30156 16454
rect 30104 16390 30156 16396
rect 30012 16244 30064 16250
rect 30012 16186 30064 16192
rect 29736 15700 29788 15706
rect 29736 15642 29788 15648
rect 30392 15570 30420 17274
rect 30484 16454 30512 17462
rect 30472 16448 30524 16454
rect 30472 16390 30524 16396
rect 30484 16114 30512 16390
rect 30472 16108 30524 16114
rect 30472 16050 30524 16056
rect 30380 15564 30432 15570
rect 30380 15506 30432 15512
rect 29736 15496 29788 15502
rect 29736 15438 29788 15444
rect 30288 15496 30340 15502
rect 30288 15438 30340 15444
rect 29552 15156 29604 15162
rect 29552 15098 29604 15104
rect 29460 15020 29512 15026
rect 29460 14962 29512 14968
rect 29184 13796 29236 13802
rect 29184 13738 29236 13744
rect 28816 13524 28868 13530
rect 28816 13466 28868 13472
rect 28816 13252 28868 13258
rect 28816 13194 28868 13200
rect 28828 12986 28856 13194
rect 29092 13184 29144 13190
rect 29092 13126 29144 13132
rect 28264 12980 28316 12986
rect 28264 12922 28316 12928
rect 28816 12980 28868 12986
rect 28816 12922 28868 12928
rect 29000 12844 29052 12850
rect 29000 12786 29052 12792
rect 28908 12368 28960 12374
rect 28908 12310 28960 12316
rect 28080 12300 28132 12306
rect 28080 12242 28132 12248
rect 27620 11756 27672 11762
rect 27620 11698 27672 11704
rect 27344 11688 27396 11694
rect 27344 11630 27396 11636
rect 27356 11286 27384 11630
rect 27344 11280 27396 11286
rect 27344 11222 27396 11228
rect 28092 11082 28120 12242
rect 28632 12164 28684 12170
rect 28632 12106 28684 12112
rect 27712 11076 27764 11082
rect 27712 11018 27764 11024
rect 28080 11076 28132 11082
rect 28080 11018 28132 11024
rect 26976 10736 27028 10742
rect 26976 10678 27028 10684
rect 26988 10606 27016 10678
rect 27068 10668 27120 10674
rect 27068 10610 27120 10616
rect 26976 10600 27028 10606
rect 26976 10542 27028 10548
rect 26424 10056 26476 10062
rect 26424 9998 26476 10004
rect 24860 9444 24912 9450
rect 24860 9386 24912 9392
rect 26252 9438 26372 9466
rect 26056 9376 26108 9382
rect 26056 9318 26108 9324
rect 24584 9036 24636 9042
rect 24584 8978 24636 8984
rect 25688 9036 25740 9042
rect 25688 8978 25740 8984
rect 24952 8900 25004 8906
rect 24952 8842 25004 8848
rect 24964 8090 24992 8842
rect 25700 8498 25728 8978
rect 26068 8974 26096 9318
rect 26252 9110 26280 9438
rect 26332 9376 26384 9382
rect 26332 9318 26384 9324
rect 26240 9104 26292 9110
rect 26240 9046 26292 9052
rect 26056 8968 26108 8974
rect 26056 8910 26108 8916
rect 25688 8492 25740 8498
rect 25688 8434 25740 8440
rect 26056 8492 26108 8498
rect 26056 8434 26108 8440
rect 24952 8084 25004 8090
rect 24952 8026 25004 8032
rect 26068 6798 26096 8434
rect 26344 7886 26372 9318
rect 26436 8634 26464 9998
rect 26424 8628 26476 8634
rect 26424 8570 26476 8576
rect 26332 7880 26384 7886
rect 26332 7822 26384 7828
rect 26056 6792 26108 6798
rect 26056 6734 26108 6740
rect 26068 5710 26096 6734
rect 26608 6316 26660 6322
rect 26608 6258 26660 6264
rect 26332 6112 26384 6118
rect 26332 6054 26384 6060
rect 26344 5778 26372 6054
rect 26332 5772 26384 5778
rect 26332 5714 26384 5720
rect 25044 5704 25096 5710
rect 25044 5646 25096 5652
rect 26056 5704 26108 5710
rect 26056 5646 26108 5652
rect 24584 3528 24636 3534
rect 24584 3470 24636 3476
rect 24596 2582 24624 3470
rect 25056 3466 25084 5646
rect 26620 5370 26648 6258
rect 26608 5364 26660 5370
rect 26608 5306 26660 5312
rect 25044 3460 25096 3466
rect 25044 3402 25096 3408
rect 24676 3392 24728 3398
rect 24676 3334 24728 3340
rect 24688 3126 24716 3334
rect 24676 3120 24728 3126
rect 24676 3062 24728 3068
rect 25056 3058 25084 3402
rect 26240 3188 26292 3194
rect 26240 3130 26292 3136
rect 25044 3052 25096 3058
rect 25044 2994 25096 3000
rect 24768 2984 24820 2990
rect 24768 2926 24820 2932
rect 24780 2650 24808 2926
rect 25228 2848 25280 2854
rect 25228 2790 25280 2796
rect 25240 2650 25268 2790
rect 24768 2644 24820 2650
rect 24768 2586 24820 2592
rect 25228 2644 25280 2650
rect 25228 2586 25280 2592
rect 24584 2576 24636 2582
rect 24584 2518 24636 2524
rect 24492 2372 24544 2378
rect 24492 2314 24544 2320
rect 26252 800 26280 3130
rect 27080 2650 27108 10610
rect 27724 10198 27752 11018
rect 28172 11008 28224 11014
rect 28172 10950 28224 10956
rect 27712 10192 27764 10198
rect 27712 10134 27764 10140
rect 27436 9988 27488 9994
rect 27436 9930 27488 9936
rect 27448 9518 27476 9930
rect 27724 9722 27752 10134
rect 28184 10062 28212 10950
rect 28644 10266 28672 12106
rect 28920 11762 28948 12310
rect 28908 11756 28960 11762
rect 28908 11698 28960 11704
rect 29012 11626 29040 12786
rect 29104 11898 29132 13126
rect 29092 11892 29144 11898
rect 29092 11834 29144 11840
rect 29000 11620 29052 11626
rect 29000 11562 29052 11568
rect 28908 11076 28960 11082
rect 28908 11018 28960 11024
rect 28816 10600 28868 10606
rect 28816 10542 28868 10548
rect 28632 10260 28684 10266
rect 28632 10202 28684 10208
rect 28172 10056 28224 10062
rect 28172 9998 28224 10004
rect 28828 9722 28856 10542
rect 27712 9716 27764 9722
rect 27712 9658 27764 9664
rect 28816 9716 28868 9722
rect 28816 9658 28868 9664
rect 27620 9648 27672 9654
rect 27620 9590 27672 9596
rect 27436 9512 27488 9518
rect 27436 9454 27488 9460
rect 27632 9178 27660 9590
rect 28920 9518 28948 11018
rect 29472 10606 29500 14962
rect 29748 14414 29776 15438
rect 29828 15360 29880 15366
rect 29828 15302 29880 15308
rect 29840 15026 29868 15302
rect 30012 15088 30064 15094
rect 30012 15030 30064 15036
rect 29828 15020 29880 15026
rect 29828 14962 29880 14968
rect 29920 14952 29972 14958
rect 29920 14894 29972 14900
rect 29932 14482 29960 14894
rect 29920 14476 29972 14482
rect 29920 14418 29972 14424
rect 30024 14414 30052 15030
rect 30300 14482 30328 15438
rect 30484 15162 30512 16050
rect 30576 15450 30604 19314
rect 31024 19304 31076 19310
rect 31024 19246 31076 19252
rect 31036 18970 31064 19246
rect 31024 18964 31076 18970
rect 31024 18906 31076 18912
rect 30748 18828 30800 18834
rect 30748 18770 30800 18776
rect 30760 16794 30788 18770
rect 30932 18080 30984 18086
rect 30932 18022 30984 18028
rect 30944 16794 30972 18022
rect 30748 16788 30800 16794
rect 30748 16730 30800 16736
rect 30932 16788 30984 16794
rect 30932 16730 30984 16736
rect 30944 16266 30972 16730
rect 30760 16238 30972 16266
rect 30760 15978 30788 16238
rect 30932 16108 30984 16114
rect 30932 16050 30984 16056
rect 30748 15972 30800 15978
rect 30748 15914 30800 15920
rect 30656 15904 30708 15910
rect 30656 15846 30708 15852
rect 30668 15570 30696 15846
rect 30656 15564 30708 15570
rect 30656 15506 30708 15512
rect 30576 15422 30696 15450
rect 30760 15434 30788 15914
rect 30472 15156 30524 15162
rect 30472 15098 30524 15104
rect 30288 14476 30340 14482
rect 30288 14418 30340 14424
rect 29736 14408 29788 14414
rect 29736 14350 29788 14356
rect 30012 14408 30064 14414
rect 30012 14350 30064 14356
rect 30300 14074 30328 14418
rect 30288 14068 30340 14074
rect 30288 14010 30340 14016
rect 30288 13932 30340 13938
rect 30288 13874 30340 13880
rect 30564 13932 30616 13938
rect 30564 13874 30616 13880
rect 30012 12776 30064 12782
rect 30012 12718 30064 12724
rect 29828 12232 29880 12238
rect 29828 12174 29880 12180
rect 29920 12232 29972 12238
rect 29920 12174 29972 12180
rect 29552 12096 29604 12102
rect 29552 12038 29604 12044
rect 29564 10742 29592 12038
rect 29840 11218 29868 12174
rect 29828 11212 29880 11218
rect 29828 11154 29880 11160
rect 29552 10736 29604 10742
rect 29552 10678 29604 10684
rect 29840 10674 29868 11154
rect 29828 10668 29880 10674
rect 29828 10610 29880 10616
rect 29460 10600 29512 10606
rect 29460 10542 29512 10548
rect 29472 10062 29500 10542
rect 29840 10130 29868 10610
rect 29932 10266 29960 12174
rect 30024 12102 30052 12718
rect 30196 12436 30248 12442
rect 30300 12434 30328 13874
rect 30472 13524 30524 13530
rect 30472 13466 30524 13472
rect 30484 12850 30512 13466
rect 30576 12986 30604 13874
rect 30564 12980 30616 12986
rect 30564 12922 30616 12928
rect 30472 12844 30524 12850
rect 30472 12786 30524 12792
rect 30248 12406 30328 12434
rect 30196 12378 30248 12384
rect 30012 12096 30064 12102
rect 30012 12038 30064 12044
rect 30024 11898 30052 12038
rect 30012 11892 30064 11898
rect 30012 11834 30064 11840
rect 30024 11354 30052 11834
rect 30104 11756 30156 11762
rect 30104 11698 30156 11704
rect 30012 11348 30064 11354
rect 30012 11290 30064 11296
rect 30116 10810 30144 11698
rect 30196 11688 30248 11694
rect 30196 11630 30248 11636
rect 30208 11286 30236 11630
rect 30196 11280 30248 11286
rect 30196 11222 30248 11228
rect 30104 10804 30156 10810
rect 30104 10746 30156 10752
rect 29920 10260 29972 10266
rect 29920 10202 29972 10208
rect 30208 10130 30236 11222
rect 30484 10810 30512 12786
rect 30668 12374 30696 15422
rect 30748 15428 30800 15434
rect 30748 15370 30800 15376
rect 30840 15360 30892 15366
rect 30840 15302 30892 15308
rect 30852 14958 30880 15302
rect 30944 15026 30972 16050
rect 30932 15020 30984 15026
rect 30932 14962 30984 14968
rect 30840 14952 30892 14958
rect 30840 14894 30892 14900
rect 31024 14272 31076 14278
rect 31024 14214 31076 14220
rect 30840 13728 30892 13734
rect 30840 13670 30892 13676
rect 30852 13190 30880 13670
rect 31036 13258 31064 14214
rect 31024 13252 31076 13258
rect 31024 13194 31076 13200
rect 30840 13184 30892 13190
rect 30840 13126 30892 13132
rect 30656 12368 30708 12374
rect 30708 12316 30788 12322
rect 30656 12310 30788 12316
rect 30668 12294 30788 12310
rect 30760 11762 30788 12294
rect 30932 12232 30984 12238
rect 30932 12174 30984 12180
rect 30748 11756 30800 11762
rect 30748 11698 30800 11704
rect 30944 11014 30972 12174
rect 30932 11008 30984 11014
rect 30932 10950 30984 10956
rect 30472 10804 30524 10810
rect 30472 10746 30524 10752
rect 30656 10668 30708 10674
rect 30656 10610 30708 10616
rect 30380 10464 30432 10470
rect 30380 10406 30432 10412
rect 29828 10124 29880 10130
rect 29828 10066 29880 10072
rect 29920 10124 29972 10130
rect 29920 10066 29972 10072
rect 30196 10124 30248 10130
rect 30196 10066 30248 10072
rect 29460 10056 29512 10062
rect 29460 9998 29512 10004
rect 29840 9586 29868 10066
rect 29828 9580 29880 9586
rect 29828 9522 29880 9528
rect 28908 9512 28960 9518
rect 28908 9454 28960 9460
rect 27620 9172 27672 9178
rect 27620 9114 27672 9120
rect 28356 9036 28408 9042
rect 28356 8978 28408 8984
rect 29184 9036 29236 9042
rect 29184 8978 29236 8984
rect 27160 8900 27212 8906
rect 27160 8842 27212 8848
rect 27620 8900 27672 8906
rect 27620 8842 27672 8848
rect 27172 8090 27200 8842
rect 27632 8634 27660 8842
rect 27620 8628 27672 8634
rect 27620 8570 27672 8576
rect 27804 8492 27856 8498
rect 27804 8434 27856 8440
rect 27988 8492 28040 8498
rect 27988 8434 28040 8440
rect 27160 8084 27212 8090
rect 27160 8026 27212 8032
rect 27344 7404 27396 7410
rect 27344 7346 27396 7352
rect 27160 7200 27212 7206
rect 27160 7142 27212 7148
rect 27172 7002 27200 7142
rect 27160 6996 27212 7002
rect 27160 6938 27212 6944
rect 27356 6458 27384 7346
rect 27816 6798 27844 8434
rect 27896 7200 27948 7206
rect 27896 7142 27948 7148
rect 27804 6792 27856 6798
rect 27804 6734 27856 6740
rect 27908 6730 27936 7142
rect 27896 6724 27948 6730
rect 27896 6666 27948 6672
rect 28000 6662 28028 8434
rect 27804 6656 27856 6662
rect 27632 6604 27804 6610
rect 27632 6598 27856 6604
rect 27988 6656 28040 6662
rect 27988 6598 28040 6604
rect 27632 6582 27844 6598
rect 27344 6452 27396 6458
rect 27344 6394 27396 6400
rect 27632 6254 27660 6582
rect 27620 6248 27672 6254
rect 27620 6190 27672 6196
rect 27632 5370 27660 6190
rect 27712 5908 27764 5914
rect 27712 5850 27764 5856
rect 27620 5364 27672 5370
rect 27620 5306 27672 5312
rect 27724 5234 27752 5850
rect 27712 5228 27764 5234
rect 27712 5170 27764 5176
rect 27528 4480 27580 4486
rect 27528 4422 27580 4428
rect 27540 4214 27568 4422
rect 27528 4208 27580 4214
rect 27528 4150 27580 4156
rect 28080 4208 28132 4214
rect 28080 4150 28132 4156
rect 27160 3936 27212 3942
rect 27160 3878 27212 3884
rect 27172 3670 27200 3878
rect 28092 3738 28120 4150
rect 28080 3732 28132 3738
rect 28080 3674 28132 3680
rect 27160 3664 27212 3670
rect 27160 3606 27212 3612
rect 28368 3534 28396 8978
rect 28632 8832 28684 8838
rect 28632 8774 28684 8780
rect 28644 8634 28672 8774
rect 28632 8628 28684 8634
rect 28632 8570 28684 8576
rect 28644 7886 28672 8570
rect 28724 8356 28776 8362
rect 28724 8298 28776 8304
rect 28632 7880 28684 7886
rect 28632 7822 28684 7828
rect 28736 7002 28764 8298
rect 28816 8288 28868 8294
rect 28816 8230 28868 8236
rect 28828 7886 28856 8230
rect 28908 7948 28960 7954
rect 28908 7890 28960 7896
rect 28816 7880 28868 7886
rect 28816 7822 28868 7828
rect 28724 6996 28776 7002
rect 28724 6938 28776 6944
rect 28736 6866 28764 6938
rect 28724 6860 28776 6866
rect 28724 6802 28776 6808
rect 28632 6792 28684 6798
rect 28920 6746 28948 7890
rect 29000 7200 29052 7206
rect 29000 7142 29052 7148
rect 28632 6734 28684 6740
rect 28448 6656 28500 6662
rect 28448 6598 28500 6604
rect 28460 6458 28488 6598
rect 28448 6452 28500 6458
rect 28448 6394 28500 6400
rect 28448 6112 28500 6118
rect 28448 6054 28500 6060
rect 28460 5710 28488 6054
rect 28448 5704 28500 5710
rect 28448 5646 28500 5652
rect 28540 5228 28592 5234
rect 28540 5170 28592 5176
rect 28448 4480 28500 4486
rect 28448 4422 28500 4428
rect 28460 4282 28488 4422
rect 28552 4282 28580 5170
rect 28644 4978 28672 6734
rect 28828 6718 28948 6746
rect 29012 6730 29040 7142
rect 29000 6724 29052 6730
rect 28828 5098 28856 6718
rect 29000 6666 29052 6672
rect 28908 6656 28960 6662
rect 28908 6598 28960 6604
rect 28920 5914 28948 6598
rect 29092 6384 29144 6390
rect 29092 6326 29144 6332
rect 29104 5914 29132 6326
rect 29196 6322 29224 8978
rect 29932 7954 29960 10066
rect 30196 9920 30248 9926
rect 30196 9862 30248 9868
rect 30208 9654 30236 9862
rect 30392 9654 30420 10406
rect 30564 10260 30616 10266
rect 30564 10202 30616 10208
rect 30196 9648 30248 9654
rect 30196 9590 30248 9596
rect 30380 9648 30432 9654
rect 30380 9590 30432 9596
rect 29920 7948 29972 7954
rect 29920 7890 29972 7896
rect 29932 6882 29960 7890
rect 30012 7472 30064 7478
rect 30012 7414 30064 7420
rect 29840 6866 29960 6882
rect 29828 6860 29960 6866
rect 29880 6854 29960 6860
rect 29828 6802 29880 6808
rect 29184 6316 29236 6322
rect 29184 6258 29236 6264
rect 28908 5908 28960 5914
rect 28908 5850 28960 5856
rect 29092 5908 29144 5914
rect 29092 5850 29144 5856
rect 29196 5710 29224 6258
rect 29840 6254 29868 6802
rect 29828 6248 29880 6254
rect 29828 6190 29880 6196
rect 30024 5914 30052 7414
rect 30104 6656 30156 6662
rect 30104 6598 30156 6604
rect 30012 5908 30064 5914
rect 30012 5850 30064 5856
rect 29736 5772 29788 5778
rect 29736 5714 29788 5720
rect 29184 5704 29236 5710
rect 29184 5646 29236 5652
rect 29644 5160 29696 5166
rect 29644 5102 29696 5108
rect 28816 5092 28868 5098
rect 28816 5034 28868 5040
rect 29000 5024 29052 5030
rect 28644 4950 28948 4978
rect 29000 4966 29052 4972
rect 29184 5024 29236 5030
rect 29184 4966 29236 4972
rect 28448 4276 28500 4282
rect 28448 4218 28500 4224
rect 28540 4276 28592 4282
rect 28540 4218 28592 4224
rect 28460 4162 28488 4218
rect 28460 4134 28580 4162
rect 28920 4146 28948 4950
rect 29012 4690 29040 4966
rect 29000 4684 29052 4690
rect 29000 4626 29052 4632
rect 29196 4622 29224 4966
rect 29184 4616 29236 4622
rect 29184 4558 29236 4564
rect 29656 4282 29684 5102
rect 29748 4622 29776 5714
rect 30116 5370 30144 6598
rect 30104 5364 30156 5370
rect 30104 5306 30156 5312
rect 30012 5092 30064 5098
rect 30012 5034 30064 5040
rect 29736 4616 29788 4622
rect 29736 4558 29788 4564
rect 29644 4276 29696 4282
rect 29644 4218 29696 4224
rect 28552 4078 28580 4134
rect 28908 4140 28960 4146
rect 28908 4082 28960 4088
rect 28540 4072 28592 4078
rect 28540 4014 28592 4020
rect 28920 3602 28948 4082
rect 29748 4010 29776 4558
rect 30024 4078 30052 5034
rect 30012 4072 30064 4078
rect 30012 4014 30064 4020
rect 29736 4004 29788 4010
rect 29736 3946 29788 3952
rect 28908 3596 28960 3602
rect 28908 3538 28960 3544
rect 28356 3528 28408 3534
rect 28356 3470 28408 3476
rect 28920 3398 28948 3538
rect 28908 3392 28960 3398
rect 28908 3334 28960 3340
rect 27068 2644 27120 2650
rect 27068 2586 27120 2592
rect 30208 2514 30236 9590
rect 30288 8560 30340 8566
rect 30288 8502 30340 8508
rect 30300 7546 30328 8502
rect 30576 8022 30604 10202
rect 30668 8634 30696 10610
rect 30840 10600 30892 10606
rect 30944 10588 30972 10950
rect 30892 10560 30972 10588
rect 30840 10542 30892 10548
rect 30852 10130 30880 10542
rect 30840 10124 30892 10130
rect 30840 10066 30892 10072
rect 30656 8628 30708 8634
rect 30656 8570 30708 8576
rect 30564 8016 30616 8022
rect 30564 7958 30616 7964
rect 30668 7954 30696 8570
rect 30852 8566 30880 10066
rect 31128 9042 31156 22918
rect 31208 21004 31260 21010
rect 31208 20946 31260 20952
rect 31220 19922 31248 20946
rect 31300 20256 31352 20262
rect 31300 20198 31352 20204
rect 31208 19916 31260 19922
rect 31208 19858 31260 19864
rect 31220 18426 31248 19858
rect 31312 19786 31340 20198
rect 31300 19780 31352 19786
rect 31300 19722 31352 19728
rect 31404 19174 31432 24618
rect 31956 24274 31984 26318
rect 32048 26042 32076 27814
rect 32036 26036 32088 26042
rect 32036 25978 32088 25984
rect 32048 24274 32076 25978
rect 31944 24268 31996 24274
rect 31944 24210 31996 24216
rect 32036 24268 32088 24274
rect 32036 24210 32088 24216
rect 31956 23662 31984 24210
rect 31944 23656 31996 23662
rect 31944 23598 31996 23604
rect 31956 23322 31984 23598
rect 32140 23526 32168 30194
rect 33060 29850 33088 30194
rect 33048 29844 33100 29850
rect 33048 29786 33100 29792
rect 32220 29640 32272 29646
rect 32220 29582 32272 29588
rect 32232 29306 32260 29582
rect 32404 29504 32456 29510
rect 32404 29446 32456 29452
rect 32220 29300 32272 29306
rect 32220 29242 32272 29248
rect 32416 28490 32444 29446
rect 33152 29306 33180 32778
rect 33324 31884 33376 31890
rect 33324 31826 33376 31832
rect 33336 30190 33364 31826
rect 33520 31362 33548 32914
rect 33612 31482 33640 34410
rect 33784 33516 33836 33522
rect 33784 33458 33836 33464
rect 33796 32434 33824 33458
rect 34532 33114 34560 37810
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 35594 37020 35902 37029
rect 35594 37018 35600 37020
rect 35656 37018 35680 37020
rect 35736 37018 35760 37020
rect 35816 37018 35840 37020
rect 35896 37018 35902 37020
rect 35656 36966 35658 37018
rect 35838 36966 35840 37018
rect 35594 36964 35600 36966
rect 35656 36964 35680 36966
rect 35736 36964 35760 36966
rect 35816 36964 35840 36966
rect 35896 36964 35902 36966
rect 35594 36955 35902 36964
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 35594 35932 35902 35941
rect 35594 35930 35600 35932
rect 35656 35930 35680 35932
rect 35736 35930 35760 35932
rect 35816 35930 35840 35932
rect 35896 35930 35902 35932
rect 35656 35878 35658 35930
rect 35838 35878 35840 35930
rect 35594 35876 35600 35878
rect 35656 35876 35680 35878
rect 35736 35876 35760 35878
rect 35816 35876 35840 35878
rect 35896 35876 35902 35878
rect 35594 35867 35902 35876
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 35594 34844 35902 34853
rect 35594 34842 35600 34844
rect 35656 34842 35680 34844
rect 35736 34842 35760 34844
rect 35816 34842 35840 34844
rect 35896 34842 35902 34844
rect 35656 34790 35658 34842
rect 35838 34790 35840 34842
rect 35594 34788 35600 34790
rect 35656 34788 35680 34790
rect 35736 34788 35760 34790
rect 35816 34788 35840 34790
rect 35896 34788 35902 34790
rect 35594 34779 35902 34788
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 35594 33756 35902 33765
rect 35594 33754 35600 33756
rect 35656 33754 35680 33756
rect 35736 33754 35760 33756
rect 35816 33754 35840 33756
rect 35896 33754 35902 33756
rect 35656 33702 35658 33754
rect 35838 33702 35840 33754
rect 35594 33700 35600 33702
rect 35656 33700 35680 33702
rect 35736 33700 35760 33702
rect 35816 33700 35840 33702
rect 35896 33700 35902 33702
rect 35594 33691 35902 33700
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 34520 33108 34572 33114
rect 34520 33050 34572 33056
rect 35594 32668 35902 32677
rect 35594 32666 35600 32668
rect 35656 32666 35680 32668
rect 35736 32666 35760 32668
rect 35816 32666 35840 32668
rect 35896 32666 35902 32668
rect 35656 32614 35658 32666
rect 35838 32614 35840 32666
rect 35594 32612 35600 32614
rect 35656 32612 35680 32614
rect 35736 32612 35760 32614
rect 35816 32612 35840 32614
rect 35896 32612 35902 32614
rect 35594 32603 35902 32612
rect 33784 32428 33836 32434
rect 33784 32370 33836 32376
rect 33692 32224 33744 32230
rect 33692 32166 33744 32172
rect 33600 31476 33652 31482
rect 33600 31418 33652 31424
rect 33520 31334 33640 31362
rect 33612 31142 33640 31334
rect 33600 31136 33652 31142
rect 33600 31078 33652 31084
rect 33612 30802 33640 31078
rect 33600 30796 33652 30802
rect 33600 30738 33652 30744
rect 33704 30666 33732 32166
rect 33796 31822 33824 32370
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 33784 31816 33836 31822
rect 33784 31758 33836 31764
rect 34520 31816 34572 31822
rect 34520 31758 34572 31764
rect 34532 31482 34560 31758
rect 35594 31580 35902 31589
rect 35594 31578 35600 31580
rect 35656 31578 35680 31580
rect 35736 31578 35760 31580
rect 35816 31578 35840 31580
rect 35896 31578 35902 31580
rect 35656 31526 35658 31578
rect 35838 31526 35840 31578
rect 35594 31524 35600 31526
rect 35656 31524 35680 31526
rect 35736 31524 35760 31526
rect 35816 31524 35840 31526
rect 35896 31524 35902 31526
rect 35594 31515 35902 31524
rect 34520 31476 34572 31482
rect 34520 31418 34572 31424
rect 34336 31340 34388 31346
rect 34336 31282 34388 31288
rect 34348 30938 34376 31282
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 34336 30932 34388 30938
rect 34336 30874 34388 30880
rect 33692 30660 33744 30666
rect 33692 30602 33744 30608
rect 33968 30592 34020 30598
rect 33968 30534 34020 30540
rect 33980 30258 34008 30534
rect 35594 30492 35902 30501
rect 35594 30490 35600 30492
rect 35656 30490 35680 30492
rect 35736 30490 35760 30492
rect 35816 30490 35840 30492
rect 35896 30490 35902 30492
rect 35656 30438 35658 30490
rect 35838 30438 35840 30490
rect 35594 30436 35600 30438
rect 35656 30436 35680 30438
rect 35736 30436 35760 30438
rect 35816 30436 35840 30438
rect 35896 30436 35902 30438
rect 35594 30427 35902 30436
rect 33968 30252 34020 30258
rect 33968 30194 34020 30200
rect 33324 30184 33376 30190
rect 33324 30126 33376 30132
rect 33980 29714 34008 30194
rect 34428 30048 34480 30054
rect 34428 29990 34480 29996
rect 33968 29708 34020 29714
rect 33968 29650 34020 29656
rect 33416 29572 33468 29578
rect 33416 29514 33468 29520
rect 33232 29504 33284 29510
rect 33232 29446 33284 29452
rect 33140 29300 33192 29306
rect 33140 29242 33192 29248
rect 32496 28960 32548 28966
rect 32496 28902 32548 28908
rect 32404 28484 32456 28490
rect 32404 28426 32456 28432
rect 32508 28150 32536 28902
rect 33152 28558 33180 29242
rect 33244 29102 33272 29446
rect 33232 29096 33284 29102
rect 33232 29038 33284 29044
rect 33244 28626 33272 29038
rect 33232 28620 33284 28626
rect 33232 28562 33284 28568
rect 33140 28552 33192 28558
rect 33140 28494 33192 28500
rect 33428 28422 33456 29514
rect 34440 29102 34468 29990
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 35594 29404 35902 29413
rect 35594 29402 35600 29404
rect 35656 29402 35680 29404
rect 35736 29402 35760 29404
rect 35816 29402 35840 29404
rect 35896 29402 35902 29404
rect 35656 29350 35658 29402
rect 35838 29350 35840 29402
rect 35594 29348 35600 29350
rect 35656 29348 35680 29350
rect 35736 29348 35760 29350
rect 35816 29348 35840 29350
rect 35896 29348 35902 29350
rect 35594 29339 35902 29348
rect 34520 29164 34572 29170
rect 34520 29106 34572 29112
rect 34428 29096 34480 29102
rect 34428 29038 34480 29044
rect 33416 28416 33468 28422
rect 33416 28358 33468 28364
rect 32496 28144 32548 28150
rect 32496 28086 32548 28092
rect 32956 28144 33008 28150
rect 32956 28086 33008 28092
rect 32508 27538 32536 28086
rect 32496 27532 32548 27538
rect 32496 27474 32548 27480
rect 32312 26988 32364 26994
rect 32312 26930 32364 26936
rect 32324 26586 32352 26930
rect 32508 26858 32536 27474
rect 32864 27464 32916 27470
rect 32864 27406 32916 27412
rect 32876 27334 32904 27406
rect 32864 27328 32916 27334
rect 32864 27270 32916 27276
rect 32496 26852 32548 26858
rect 32496 26794 32548 26800
rect 32312 26580 32364 26586
rect 32312 26522 32364 26528
rect 32324 25786 32352 26522
rect 32588 26308 32640 26314
rect 32588 26250 32640 26256
rect 32600 25906 32628 26250
rect 32876 26234 32904 27270
rect 32968 27130 32996 28086
rect 33324 27940 33376 27946
rect 33324 27882 33376 27888
rect 33336 27538 33364 27882
rect 33324 27532 33376 27538
rect 33324 27474 33376 27480
rect 33048 27396 33100 27402
rect 33048 27338 33100 27344
rect 32956 27124 33008 27130
rect 32956 27066 33008 27072
rect 32968 26926 32996 27066
rect 32956 26920 33008 26926
rect 32956 26862 33008 26868
rect 32956 26784 33008 26790
rect 32956 26726 33008 26732
rect 32968 26382 32996 26726
rect 33060 26450 33088 27338
rect 33336 27146 33364 27474
rect 33152 27130 33364 27146
rect 33152 27124 33376 27130
rect 33152 27118 33324 27124
rect 33048 26444 33100 26450
rect 33048 26386 33100 26392
rect 33152 26382 33180 27118
rect 33324 27066 33376 27072
rect 33336 27035 33364 27066
rect 33428 26518 33456 28358
rect 33508 28212 33560 28218
rect 33508 28154 33560 28160
rect 33520 27062 33548 28154
rect 34440 28150 34468 29038
rect 34532 28762 34560 29106
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34520 28756 34572 28762
rect 34520 28698 34572 28704
rect 35072 28552 35124 28558
rect 35072 28494 35124 28500
rect 35440 28552 35492 28558
rect 35440 28494 35492 28500
rect 34612 28416 34664 28422
rect 34612 28358 34664 28364
rect 34428 28144 34480 28150
rect 34428 28086 34480 28092
rect 34440 27690 34468 28086
rect 34440 27662 34560 27690
rect 33508 27056 33560 27062
rect 33508 26998 33560 27004
rect 34244 26988 34296 26994
rect 34244 26930 34296 26936
rect 33968 26784 34020 26790
rect 33968 26726 34020 26732
rect 33416 26512 33468 26518
rect 33416 26454 33468 26460
rect 32956 26376 33008 26382
rect 32956 26318 33008 26324
rect 33140 26376 33192 26382
rect 33140 26318 33192 26324
rect 33428 26234 33456 26454
rect 33876 26444 33928 26450
rect 33876 26386 33928 26392
rect 32876 26206 33088 26234
rect 33060 25974 33088 26206
rect 33336 26206 33456 26234
rect 33692 26240 33744 26246
rect 33048 25968 33100 25974
rect 33048 25910 33100 25916
rect 32588 25900 32640 25906
rect 32588 25842 32640 25848
rect 32324 25770 32444 25786
rect 32324 25764 32456 25770
rect 32324 25758 32404 25764
rect 32324 25226 32352 25758
rect 32404 25706 32456 25712
rect 32600 25498 32628 25842
rect 32772 25696 32824 25702
rect 32772 25638 32824 25644
rect 32588 25492 32640 25498
rect 32588 25434 32640 25440
rect 32312 25220 32364 25226
rect 32312 25162 32364 25168
rect 32496 24812 32548 24818
rect 32496 24754 32548 24760
rect 32220 24744 32272 24750
rect 32220 24686 32272 24692
rect 32232 24206 32260 24686
rect 32508 24274 32536 24754
rect 32312 24268 32364 24274
rect 32312 24210 32364 24216
rect 32496 24268 32548 24274
rect 32496 24210 32548 24216
rect 32220 24200 32272 24206
rect 32220 24142 32272 24148
rect 32128 23520 32180 23526
rect 32128 23462 32180 23468
rect 31944 23316 31996 23322
rect 31944 23258 31996 23264
rect 32232 23050 32260 24142
rect 32324 23644 32352 24210
rect 32508 23730 32536 24210
rect 32496 23724 32548 23730
rect 32496 23666 32548 23672
rect 32404 23656 32456 23662
rect 32324 23616 32404 23644
rect 32404 23598 32456 23604
rect 32312 23520 32364 23526
rect 32312 23462 32364 23468
rect 32220 23044 32272 23050
rect 32220 22986 32272 22992
rect 31760 22704 31812 22710
rect 31760 22646 31812 22652
rect 31772 22098 31800 22646
rect 31944 22228 31996 22234
rect 31944 22170 31996 22176
rect 31760 22092 31812 22098
rect 31760 22034 31812 22040
rect 31956 22030 31984 22170
rect 31944 22024 31996 22030
rect 31944 21966 31996 21972
rect 31484 21412 31536 21418
rect 31484 21354 31536 21360
rect 31496 21078 31524 21354
rect 31484 21072 31536 21078
rect 31484 21014 31536 21020
rect 31576 20936 31628 20942
rect 31576 20878 31628 20884
rect 31588 20602 31616 20878
rect 31576 20596 31628 20602
rect 31576 20538 31628 20544
rect 31576 20460 31628 20466
rect 31576 20402 31628 20408
rect 31588 19378 31616 20402
rect 31576 19372 31628 19378
rect 31576 19314 31628 19320
rect 31392 19168 31444 19174
rect 31392 19110 31444 19116
rect 31852 19168 31904 19174
rect 31852 19110 31904 19116
rect 31864 18766 31892 19110
rect 32324 18766 32352 23462
rect 32416 22098 32444 23598
rect 32508 23186 32536 23666
rect 32784 23322 32812 25638
rect 33060 25294 33088 25910
rect 33336 25906 33364 26206
rect 33692 26182 33744 26188
rect 33140 25900 33192 25906
rect 33140 25842 33192 25848
rect 33324 25900 33376 25906
rect 33324 25842 33376 25848
rect 33048 25288 33100 25294
rect 33048 25230 33100 25236
rect 33152 24206 33180 25842
rect 33704 25226 33732 26182
rect 33888 26042 33916 26386
rect 33980 26382 34008 26726
rect 34256 26586 34284 26930
rect 34244 26580 34296 26586
rect 34244 26522 34296 26528
rect 34532 26450 34560 27662
rect 34624 27606 34652 28358
rect 35084 28218 35112 28494
rect 35164 28416 35216 28422
rect 35164 28358 35216 28364
rect 35072 28212 35124 28218
rect 35072 28154 35124 28160
rect 35176 28150 35204 28358
rect 35164 28144 35216 28150
rect 35164 28086 35216 28092
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 35452 27674 35480 28494
rect 35594 28316 35902 28325
rect 35594 28314 35600 28316
rect 35656 28314 35680 28316
rect 35736 28314 35760 28316
rect 35816 28314 35840 28316
rect 35896 28314 35902 28316
rect 35656 28262 35658 28314
rect 35838 28262 35840 28314
rect 35594 28260 35600 28262
rect 35656 28260 35680 28262
rect 35736 28260 35760 28262
rect 35816 28260 35840 28262
rect 35896 28260 35902 28262
rect 35594 28251 35902 28260
rect 35440 27668 35492 27674
rect 35440 27610 35492 27616
rect 34612 27600 34664 27606
rect 34612 27542 34664 27548
rect 34796 27532 34848 27538
rect 34796 27474 34848 27480
rect 35164 27532 35216 27538
rect 35164 27474 35216 27480
rect 34808 26926 34836 27474
rect 35176 27334 35204 27474
rect 35164 27328 35216 27334
rect 35164 27270 35216 27276
rect 35594 27228 35902 27237
rect 35594 27226 35600 27228
rect 35656 27226 35680 27228
rect 35736 27226 35760 27228
rect 35816 27226 35840 27228
rect 35896 27226 35902 27228
rect 35656 27174 35658 27226
rect 35838 27174 35840 27226
rect 35594 27172 35600 27174
rect 35656 27172 35680 27174
rect 35736 27172 35760 27174
rect 35816 27172 35840 27174
rect 35896 27172 35902 27174
rect 35594 27163 35902 27172
rect 35808 26988 35860 26994
rect 35808 26930 35860 26936
rect 34796 26920 34848 26926
rect 34796 26862 34848 26868
rect 34612 26852 34664 26858
rect 34612 26794 34664 26800
rect 34704 26852 34756 26858
rect 34704 26794 34756 26800
rect 34624 26518 34652 26794
rect 34612 26512 34664 26518
rect 34612 26454 34664 26460
rect 34520 26444 34572 26450
rect 34520 26386 34572 26392
rect 33968 26376 34020 26382
rect 34716 26330 34744 26794
rect 34808 26790 34836 26862
rect 34796 26784 34848 26790
rect 34796 26726 34848 26732
rect 35440 26784 35492 26790
rect 35440 26726 35492 26732
rect 35624 26784 35676 26790
rect 35624 26726 35676 26732
rect 33968 26318 34020 26324
rect 34520 26308 34572 26314
rect 34520 26250 34572 26256
rect 34624 26302 34744 26330
rect 33876 26036 33928 26042
rect 33876 25978 33928 25984
rect 34532 25770 34560 26250
rect 34624 25906 34652 26302
rect 34808 26234 34836 26726
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 35348 26376 35400 26382
rect 35348 26318 35400 26324
rect 34716 26206 34836 26234
rect 34612 25900 34664 25906
rect 34612 25842 34664 25848
rect 34716 25786 34744 26206
rect 34520 25764 34572 25770
rect 34520 25706 34572 25712
rect 34624 25758 34744 25786
rect 35360 25786 35388 26318
rect 35452 25888 35480 26726
rect 35636 26450 35664 26726
rect 35820 26586 35848 26930
rect 35808 26580 35860 26586
rect 35808 26522 35860 26528
rect 35624 26444 35676 26450
rect 35624 26386 35676 26392
rect 35594 26140 35902 26149
rect 35594 26138 35600 26140
rect 35656 26138 35680 26140
rect 35736 26138 35760 26140
rect 35816 26138 35840 26140
rect 35896 26138 35902 26140
rect 35656 26086 35658 26138
rect 35838 26086 35840 26138
rect 35594 26084 35600 26086
rect 35656 26084 35680 26086
rect 35736 26084 35760 26086
rect 35816 26084 35840 26086
rect 35896 26084 35902 26086
rect 35594 26075 35902 26084
rect 35452 25860 35572 25888
rect 35360 25758 35480 25786
rect 34244 25288 34296 25294
rect 34244 25230 34296 25236
rect 33232 25220 33284 25226
rect 33232 25162 33284 25168
rect 33692 25220 33744 25226
rect 33692 25162 33744 25168
rect 34152 25220 34204 25226
rect 34152 25162 34204 25168
rect 33244 24818 33272 25162
rect 33232 24812 33284 24818
rect 33232 24754 33284 24760
rect 33140 24200 33192 24206
rect 33140 24142 33192 24148
rect 32772 23316 32824 23322
rect 32772 23258 32824 23264
rect 32496 23180 32548 23186
rect 32496 23122 32548 23128
rect 32784 22710 32812 23258
rect 32956 23044 33008 23050
rect 32956 22986 33008 22992
rect 32968 22710 32996 22986
rect 33152 22778 33180 24142
rect 33244 23866 33272 24754
rect 33508 24744 33560 24750
rect 33508 24686 33560 24692
rect 33520 24342 33548 24686
rect 33508 24336 33560 24342
rect 33508 24278 33560 24284
rect 33232 23860 33284 23866
rect 33232 23802 33284 23808
rect 33520 23730 33548 24278
rect 33600 24064 33652 24070
rect 33600 24006 33652 24012
rect 33508 23724 33560 23730
rect 33508 23666 33560 23672
rect 33612 23662 33640 24006
rect 33600 23656 33652 23662
rect 33600 23598 33652 23604
rect 33508 23316 33560 23322
rect 33508 23258 33560 23264
rect 33140 22772 33192 22778
rect 33140 22714 33192 22720
rect 32772 22704 32824 22710
rect 32772 22646 32824 22652
rect 32956 22704 33008 22710
rect 32956 22646 33008 22652
rect 32588 22228 32640 22234
rect 32588 22170 32640 22176
rect 32404 22092 32456 22098
rect 32404 22034 32456 22040
rect 32416 21486 32444 22034
rect 32600 21554 32628 22170
rect 32864 21956 32916 21962
rect 32864 21898 32916 21904
rect 32876 21690 32904 21898
rect 32864 21684 32916 21690
rect 32864 21626 32916 21632
rect 32496 21548 32548 21554
rect 32496 21490 32548 21496
rect 32588 21548 32640 21554
rect 32588 21490 32640 21496
rect 32404 21480 32456 21486
rect 32404 21422 32456 21428
rect 32416 21146 32444 21422
rect 32404 21140 32456 21146
rect 32404 21082 32456 21088
rect 32508 20058 32536 21490
rect 32876 20942 32904 21626
rect 32864 20936 32916 20942
rect 32864 20878 32916 20884
rect 32876 20466 32904 20878
rect 32864 20460 32916 20466
rect 32864 20402 32916 20408
rect 32496 20052 32548 20058
rect 32496 19994 32548 20000
rect 32772 19440 32824 19446
rect 32772 19382 32824 19388
rect 32784 18970 32812 19382
rect 32772 18964 32824 18970
rect 32772 18906 32824 18912
rect 31852 18760 31904 18766
rect 31852 18702 31904 18708
rect 32312 18760 32364 18766
rect 32312 18702 32364 18708
rect 31300 18692 31352 18698
rect 31300 18634 31352 18640
rect 31208 18420 31260 18426
rect 31208 18362 31260 18368
rect 31220 17746 31248 18362
rect 31312 18154 31340 18634
rect 31760 18420 31812 18426
rect 31760 18362 31812 18368
rect 32404 18420 32456 18426
rect 32404 18362 32456 18368
rect 31300 18148 31352 18154
rect 31300 18090 31352 18096
rect 31772 18086 31800 18362
rect 31760 18080 31812 18086
rect 31760 18022 31812 18028
rect 31208 17740 31260 17746
rect 31208 17682 31260 17688
rect 31220 17338 31248 17682
rect 31208 17332 31260 17338
rect 31208 17274 31260 17280
rect 31668 17264 31720 17270
rect 31668 17206 31720 17212
rect 31680 16590 31708 17206
rect 32416 16998 32444 18362
rect 32680 17740 32732 17746
rect 32680 17682 32732 17688
rect 31852 16992 31904 16998
rect 31852 16934 31904 16940
rect 32404 16992 32456 16998
rect 32404 16934 32456 16940
rect 31668 16584 31720 16590
rect 31668 16526 31720 16532
rect 31864 16522 31892 16934
rect 32692 16590 32720 17682
rect 32968 17678 32996 22646
rect 33152 22574 33180 22714
rect 33140 22568 33192 22574
rect 33140 22510 33192 22516
rect 33152 21962 33180 22510
rect 33520 22234 33548 23258
rect 33600 23112 33652 23118
rect 33600 23054 33652 23060
rect 33508 22228 33560 22234
rect 33508 22170 33560 22176
rect 33140 21956 33192 21962
rect 33140 21898 33192 21904
rect 33416 21888 33468 21894
rect 33416 21830 33468 21836
rect 33428 20874 33456 21830
rect 33520 21622 33548 22170
rect 33612 22166 33640 23054
rect 33704 22642 33732 25162
rect 33784 24608 33836 24614
rect 33784 24550 33836 24556
rect 33968 24608 34020 24614
rect 33968 24550 34020 24556
rect 33796 23118 33824 24550
rect 33784 23112 33836 23118
rect 33784 23054 33836 23060
rect 33692 22636 33744 22642
rect 33692 22578 33744 22584
rect 33600 22160 33652 22166
rect 33600 22102 33652 22108
rect 33704 22098 33732 22578
rect 33692 22092 33744 22098
rect 33692 22034 33744 22040
rect 33600 22024 33652 22030
rect 33796 21978 33824 23054
rect 33980 22506 34008 24550
rect 34164 24274 34192 25162
rect 34256 25158 34284 25230
rect 34244 25152 34296 25158
rect 34244 25094 34296 25100
rect 34624 24682 34652 25758
rect 35452 25702 35480 25758
rect 35440 25696 35492 25702
rect 35440 25638 35492 25644
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 34796 25152 34848 25158
rect 34796 25094 34848 25100
rect 34808 24954 34836 25094
rect 34796 24948 34848 24954
rect 34796 24890 34848 24896
rect 34704 24744 34756 24750
rect 34704 24686 34756 24692
rect 34612 24676 34664 24682
rect 34612 24618 34664 24624
rect 34624 24274 34652 24618
rect 34716 24342 34744 24686
rect 35348 24608 35400 24614
rect 35348 24550 35400 24556
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 34704 24336 34756 24342
rect 34704 24278 34756 24284
rect 34152 24268 34204 24274
rect 34152 24210 34204 24216
rect 34612 24268 34664 24274
rect 34612 24210 34664 24216
rect 34428 24064 34480 24070
rect 34428 24006 34480 24012
rect 34440 23730 34468 24006
rect 34428 23724 34480 23730
rect 34428 23666 34480 23672
rect 33968 22500 34020 22506
rect 33968 22442 34020 22448
rect 33980 22030 34008 22442
rect 34428 22228 34480 22234
rect 34428 22170 34480 22176
rect 34440 22098 34468 22170
rect 34428 22092 34480 22098
rect 34428 22034 34480 22040
rect 33652 21972 33824 21978
rect 33600 21966 33824 21972
rect 33968 22024 34020 22030
rect 33968 21966 34020 21972
rect 33612 21950 33824 21966
rect 33600 21888 33652 21894
rect 33600 21830 33652 21836
rect 33508 21616 33560 21622
rect 33508 21558 33560 21564
rect 33520 20874 33548 21558
rect 33612 20942 33640 21830
rect 33692 21480 33744 21486
rect 33692 21422 33744 21428
rect 34336 21480 34388 21486
rect 34336 21422 34388 21428
rect 33704 21146 33732 21422
rect 34060 21344 34112 21350
rect 34060 21286 34112 21292
rect 33692 21140 33744 21146
rect 33692 21082 33744 21088
rect 34072 20942 34100 21286
rect 33600 20936 33652 20942
rect 33600 20878 33652 20884
rect 34060 20936 34112 20942
rect 34060 20878 34112 20884
rect 33416 20868 33468 20874
rect 33416 20810 33468 20816
rect 33508 20868 33560 20874
rect 33508 20810 33560 20816
rect 33428 20398 33456 20810
rect 33784 20800 33836 20806
rect 33784 20742 33836 20748
rect 34152 20800 34204 20806
rect 34152 20742 34204 20748
rect 33796 20398 33824 20742
rect 34164 20466 34192 20742
rect 34152 20460 34204 20466
rect 34152 20402 34204 20408
rect 33416 20392 33468 20398
rect 33416 20334 33468 20340
rect 33784 20392 33836 20398
rect 33784 20334 33836 20340
rect 34060 20256 34112 20262
rect 34060 20198 34112 20204
rect 34072 19922 34100 20198
rect 34348 19922 34376 21422
rect 34624 21078 34652 24210
rect 34716 23322 34744 24278
rect 34980 24064 35032 24070
rect 34980 24006 35032 24012
rect 34992 23730 35020 24006
rect 34980 23724 35032 23730
rect 34980 23666 35032 23672
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 34704 23316 34756 23322
rect 34704 23258 34756 23264
rect 35360 23202 35388 24550
rect 35452 23798 35480 25638
rect 35544 25294 35572 25860
rect 35532 25288 35584 25294
rect 35532 25230 35584 25236
rect 35594 25052 35902 25061
rect 35594 25050 35600 25052
rect 35656 25050 35680 25052
rect 35736 25050 35760 25052
rect 35816 25050 35840 25052
rect 35896 25050 35902 25052
rect 35656 24998 35658 25050
rect 35838 24998 35840 25050
rect 35594 24996 35600 24998
rect 35656 24996 35680 24998
rect 35736 24996 35760 24998
rect 35816 24996 35840 24998
rect 35896 24996 35902 24998
rect 35594 24987 35902 24996
rect 35594 23964 35902 23973
rect 35594 23962 35600 23964
rect 35656 23962 35680 23964
rect 35736 23962 35760 23964
rect 35816 23962 35840 23964
rect 35896 23962 35902 23964
rect 35656 23910 35658 23962
rect 35838 23910 35840 23962
rect 35594 23908 35600 23910
rect 35656 23908 35680 23910
rect 35736 23908 35760 23910
rect 35816 23908 35840 23910
rect 35896 23908 35902 23910
rect 35594 23899 35902 23908
rect 35440 23792 35492 23798
rect 35440 23734 35492 23740
rect 35268 23174 35388 23202
rect 35452 23186 35480 23734
rect 35440 23180 35492 23186
rect 35268 22574 35296 23174
rect 35440 23122 35492 23128
rect 35348 23044 35400 23050
rect 35348 22986 35400 22992
rect 35256 22568 35308 22574
rect 35256 22510 35308 22516
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 34796 22160 34848 22166
rect 34796 22102 34848 22108
rect 34808 21350 34836 22102
rect 35360 22098 35388 22986
rect 35992 22976 36044 22982
rect 35992 22918 36044 22924
rect 35594 22876 35902 22885
rect 35594 22874 35600 22876
rect 35656 22874 35680 22876
rect 35736 22874 35760 22876
rect 35816 22874 35840 22876
rect 35896 22874 35902 22876
rect 35656 22822 35658 22874
rect 35838 22822 35840 22874
rect 35594 22820 35600 22822
rect 35656 22820 35680 22822
rect 35736 22820 35760 22822
rect 35816 22820 35840 22822
rect 35896 22820 35902 22822
rect 35594 22811 35902 22820
rect 36004 22778 36032 22918
rect 35992 22772 36044 22778
rect 35992 22714 36044 22720
rect 36096 22710 36124 40174
rect 37002 40093 37058 40174
rect 36910 38720 36966 38729
rect 36910 38655 36966 38664
rect 36924 38554 36952 38655
rect 36912 38548 36964 38554
rect 36912 38490 36964 38496
rect 36912 35080 36964 35086
rect 36912 35022 36964 35028
rect 37094 35048 37150 35057
rect 36924 31482 36952 35022
rect 37094 34983 37150 34992
rect 37108 34950 37136 34983
rect 37096 34944 37148 34950
rect 37096 34886 37148 34892
rect 37096 31680 37148 31686
rect 37096 31622 37148 31628
rect 36912 31476 36964 31482
rect 36912 31418 36964 31424
rect 37108 31385 37136 31622
rect 37094 31376 37150 31385
rect 37094 31311 37150 31320
rect 36176 28144 36228 28150
rect 36176 28086 36228 28092
rect 36188 27606 36216 28086
rect 36636 27872 36688 27878
rect 36636 27814 36688 27820
rect 36176 27600 36228 27606
rect 36176 27542 36228 27548
rect 36648 27538 36676 27814
rect 37094 27704 37150 27713
rect 37094 27639 37150 27648
rect 37108 27606 37136 27639
rect 37096 27600 37148 27606
rect 37096 27542 37148 27548
rect 36636 27532 36688 27538
rect 36636 27474 36688 27480
rect 36360 27464 36412 27470
rect 36360 27406 36412 27412
rect 37004 27464 37056 27470
rect 37004 27406 37056 27412
rect 36268 25968 36320 25974
rect 36268 25910 36320 25916
rect 36176 25832 36228 25838
rect 36176 25774 36228 25780
rect 36188 25498 36216 25774
rect 36280 25498 36308 25910
rect 36176 25492 36228 25498
rect 36176 25434 36228 25440
rect 36268 25492 36320 25498
rect 36268 25434 36320 25440
rect 36372 25294 36400 27406
rect 36452 27328 36504 27334
rect 36452 27270 36504 27276
rect 36464 26994 36492 27270
rect 36452 26988 36504 26994
rect 36452 26930 36504 26936
rect 36452 26308 36504 26314
rect 36452 26250 36504 26256
rect 36360 25288 36412 25294
rect 36360 25230 36412 25236
rect 36372 24818 36400 25230
rect 36464 24818 36492 26250
rect 36360 24812 36412 24818
rect 36360 24754 36412 24760
rect 36452 24812 36504 24818
rect 36452 24754 36504 24760
rect 36912 24200 36964 24206
rect 36912 24142 36964 24148
rect 36820 24132 36872 24138
rect 36820 24074 36872 24080
rect 36832 23866 36860 24074
rect 36820 23860 36872 23866
rect 36820 23802 36872 23808
rect 36452 23724 36504 23730
rect 36452 23666 36504 23672
rect 36464 22778 36492 23666
rect 36452 22772 36504 22778
rect 36452 22714 36504 22720
rect 36084 22704 36136 22710
rect 36084 22646 36136 22652
rect 36544 22636 36596 22642
rect 36544 22578 36596 22584
rect 35348 22092 35400 22098
rect 35348 22034 35400 22040
rect 36556 22030 36584 22578
rect 36924 22094 36952 24142
rect 36832 22066 36952 22094
rect 36084 22024 36136 22030
rect 36084 21966 36136 21972
rect 36544 22024 36596 22030
rect 36544 21966 36596 21972
rect 35992 21888 36044 21894
rect 35992 21830 36044 21836
rect 35594 21788 35902 21797
rect 35594 21786 35600 21788
rect 35656 21786 35680 21788
rect 35736 21786 35760 21788
rect 35816 21786 35840 21788
rect 35896 21786 35902 21788
rect 35656 21734 35658 21786
rect 35838 21734 35840 21786
rect 35594 21732 35600 21734
rect 35656 21732 35680 21734
rect 35736 21732 35760 21734
rect 35816 21732 35840 21734
rect 35896 21732 35902 21734
rect 35594 21723 35902 21732
rect 36004 21622 36032 21830
rect 35992 21616 36044 21622
rect 35992 21558 36044 21564
rect 35348 21480 35400 21486
rect 35348 21422 35400 21428
rect 34796 21344 34848 21350
rect 34796 21286 34848 21292
rect 34612 21072 34664 21078
rect 34612 21014 34664 21020
rect 34808 21010 34836 21286
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34796 21004 34848 21010
rect 34796 20946 34848 20952
rect 34980 20800 35032 20806
rect 34980 20742 35032 20748
rect 34992 20466 35020 20742
rect 35360 20602 35388 21422
rect 35594 20700 35902 20709
rect 35594 20698 35600 20700
rect 35656 20698 35680 20700
rect 35736 20698 35760 20700
rect 35816 20698 35840 20700
rect 35896 20698 35902 20700
rect 35656 20646 35658 20698
rect 35838 20646 35840 20698
rect 35594 20644 35600 20646
rect 35656 20644 35680 20646
rect 35736 20644 35760 20646
rect 35816 20644 35840 20646
rect 35896 20644 35902 20646
rect 35594 20635 35902 20644
rect 35348 20596 35400 20602
rect 35348 20538 35400 20544
rect 36096 20534 36124 21966
rect 36084 20528 36136 20534
rect 36084 20470 36136 20476
rect 34980 20460 35032 20466
rect 34980 20402 35032 20408
rect 36636 20460 36688 20466
rect 36636 20402 36688 20408
rect 35716 20256 35768 20262
rect 35716 20198 35768 20204
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 34060 19916 34112 19922
rect 34060 19858 34112 19864
rect 34336 19916 34388 19922
rect 34336 19858 34388 19864
rect 34348 19378 34376 19858
rect 35728 19786 35756 20198
rect 35716 19780 35768 19786
rect 35716 19722 35768 19728
rect 35594 19612 35902 19621
rect 35594 19610 35600 19612
rect 35656 19610 35680 19612
rect 35736 19610 35760 19612
rect 35816 19610 35840 19612
rect 35896 19610 35902 19612
rect 35656 19558 35658 19610
rect 35838 19558 35840 19610
rect 35594 19556 35600 19558
rect 35656 19556 35680 19558
rect 35736 19556 35760 19558
rect 35816 19556 35840 19558
rect 35896 19556 35902 19558
rect 35594 19547 35902 19556
rect 34336 19372 34388 19378
rect 34336 19314 34388 19320
rect 33416 18760 33468 18766
rect 33416 18702 33468 18708
rect 33428 18290 33456 18702
rect 34348 18358 34376 19314
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 35072 18624 35124 18630
rect 35072 18566 35124 18572
rect 35084 18358 35112 18566
rect 35594 18524 35902 18533
rect 35594 18522 35600 18524
rect 35656 18522 35680 18524
rect 35736 18522 35760 18524
rect 35816 18522 35840 18524
rect 35896 18522 35902 18524
rect 35656 18470 35658 18522
rect 35838 18470 35840 18522
rect 35594 18468 35600 18470
rect 35656 18468 35680 18470
rect 35736 18468 35760 18470
rect 35816 18468 35840 18470
rect 35896 18468 35902 18470
rect 35594 18459 35902 18468
rect 34336 18352 34388 18358
rect 34336 18294 34388 18300
rect 35072 18352 35124 18358
rect 35072 18294 35124 18300
rect 33416 18284 33468 18290
rect 33416 18226 33468 18232
rect 32956 17672 33008 17678
rect 32956 17614 33008 17620
rect 33232 17264 33284 17270
rect 33232 17206 33284 17212
rect 33244 16590 33272 17206
rect 33324 17128 33376 17134
rect 33324 17070 33376 17076
rect 32680 16584 32732 16590
rect 32680 16526 32732 16532
rect 33232 16584 33284 16590
rect 33232 16526 33284 16532
rect 31852 16516 31904 16522
rect 31852 16458 31904 16464
rect 33336 16454 33364 17070
rect 33428 16658 33456 18226
rect 34060 18216 34112 18222
rect 34060 18158 34112 18164
rect 34072 17882 34100 18158
rect 34060 17876 34112 17882
rect 34060 17818 34112 17824
rect 34060 17672 34112 17678
rect 34060 17614 34112 17620
rect 34072 17134 34100 17614
rect 34348 17338 34376 18294
rect 34796 18080 34848 18086
rect 34796 18022 34848 18028
rect 34808 17746 34836 18022
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 34796 17740 34848 17746
rect 34796 17682 34848 17688
rect 34336 17332 34388 17338
rect 34336 17274 34388 17280
rect 34348 17202 34376 17274
rect 34336 17196 34388 17202
rect 34336 17138 34388 17144
rect 34060 17128 34112 17134
rect 34060 17070 34112 17076
rect 34072 16658 34100 17070
rect 33416 16652 33468 16658
rect 33416 16594 33468 16600
rect 34060 16652 34112 16658
rect 34060 16594 34112 16600
rect 33324 16448 33376 16454
rect 33324 16390 33376 16396
rect 32772 16176 32824 16182
rect 32772 16118 32824 16124
rect 31484 16108 31536 16114
rect 31484 16050 31536 16056
rect 32496 16108 32548 16114
rect 32496 16050 32548 16056
rect 32680 16108 32732 16114
rect 32680 16050 32732 16056
rect 31496 15366 31524 16050
rect 32404 15904 32456 15910
rect 32404 15846 32456 15852
rect 31760 15496 31812 15502
rect 31760 15438 31812 15444
rect 31484 15360 31536 15366
rect 31484 15302 31536 15308
rect 31576 14884 31628 14890
rect 31576 14826 31628 14832
rect 31208 14816 31260 14822
rect 31208 14758 31260 14764
rect 31220 14550 31248 14758
rect 31208 14544 31260 14550
rect 31208 14486 31260 14492
rect 31588 14482 31616 14826
rect 31772 14618 31800 15438
rect 32128 15088 32180 15094
rect 32128 15030 32180 15036
rect 32140 14822 32168 15030
rect 32128 14816 32180 14822
rect 32128 14758 32180 14764
rect 31760 14612 31812 14618
rect 31760 14554 31812 14560
rect 31576 14476 31628 14482
rect 31576 14418 31628 14424
rect 32416 14414 32444 15846
rect 32508 15706 32536 16050
rect 32496 15700 32548 15706
rect 32496 15642 32548 15648
rect 32508 14958 32536 15642
rect 32692 15178 32720 16050
rect 32784 15366 32812 16118
rect 33336 15706 33364 16390
rect 33324 15700 33376 15706
rect 33324 15642 33376 15648
rect 33428 15586 33456 16594
rect 33336 15558 33456 15586
rect 34348 15570 34376 17138
rect 34808 16794 34836 17682
rect 35072 17604 35124 17610
rect 35072 17546 35124 17552
rect 35348 17604 35400 17610
rect 35348 17546 35400 17552
rect 35084 17338 35112 17546
rect 35256 17536 35308 17542
rect 35256 17478 35308 17484
rect 35072 17332 35124 17338
rect 35072 17274 35124 17280
rect 35268 17270 35296 17478
rect 35256 17264 35308 17270
rect 35256 17206 35308 17212
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 35360 16794 35388 17546
rect 35594 17436 35902 17445
rect 35594 17434 35600 17436
rect 35656 17434 35680 17436
rect 35736 17434 35760 17436
rect 35816 17434 35840 17436
rect 35896 17434 35902 17436
rect 35656 17382 35658 17434
rect 35838 17382 35840 17434
rect 35594 17380 35600 17382
rect 35656 17380 35680 17382
rect 35736 17380 35760 17382
rect 35816 17380 35840 17382
rect 35896 17380 35902 17382
rect 35594 17371 35902 17380
rect 35440 17332 35492 17338
rect 35440 17274 35492 17280
rect 34796 16788 34848 16794
rect 34796 16730 34848 16736
rect 35348 16788 35400 16794
rect 35348 16730 35400 16736
rect 35360 16114 35388 16730
rect 35452 16522 35480 17274
rect 35900 17264 35952 17270
rect 35900 17206 35952 17212
rect 35912 16794 35940 17206
rect 35900 16788 35952 16794
rect 35900 16730 35952 16736
rect 36176 16584 36228 16590
rect 36176 16526 36228 16532
rect 35440 16516 35492 16522
rect 35440 16458 35492 16464
rect 35452 16182 35480 16458
rect 35594 16348 35902 16357
rect 35594 16346 35600 16348
rect 35656 16346 35680 16348
rect 35736 16346 35760 16348
rect 35816 16346 35840 16348
rect 35896 16346 35902 16348
rect 35656 16294 35658 16346
rect 35838 16294 35840 16346
rect 35594 16292 35600 16294
rect 35656 16292 35680 16294
rect 35736 16292 35760 16294
rect 35816 16292 35840 16294
rect 35896 16292 35902 16294
rect 35594 16283 35902 16292
rect 35440 16176 35492 16182
rect 35440 16118 35492 16124
rect 36188 16114 36216 16526
rect 35348 16108 35400 16114
rect 35348 16050 35400 16056
rect 36176 16108 36228 16114
rect 36176 16050 36228 16056
rect 34520 16040 34572 16046
rect 34520 15982 34572 15988
rect 34336 15564 34388 15570
rect 33048 15428 33100 15434
rect 33048 15370 33100 15376
rect 32772 15360 32824 15366
rect 32772 15302 32824 15308
rect 32600 15162 32720 15178
rect 32588 15156 32720 15162
rect 32640 15150 32720 15156
rect 32588 15098 32640 15104
rect 32496 14952 32548 14958
rect 32496 14894 32548 14900
rect 32508 14822 32536 14894
rect 32496 14816 32548 14822
rect 32496 14758 32548 14764
rect 32692 14482 32720 15150
rect 32784 15094 32812 15302
rect 33060 15162 33088 15370
rect 33048 15156 33100 15162
rect 33048 15098 33100 15104
rect 32772 15088 32824 15094
rect 32772 15030 32824 15036
rect 33336 15026 33364 15558
rect 34336 15506 34388 15512
rect 34060 15428 34112 15434
rect 34060 15370 34112 15376
rect 33324 15020 33376 15026
rect 33324 14962 33376 14968
rect 32680 14476 32732 14482
rect 32680 14418 32732 14424
rect 31392 14408 31444 14414
rect 31392 14350 31444 14356
rect 32404 14408 32456 14414
rect 32404 14350 32456 14356
rect 33232 14408 33284 14414
rect 33232 14350 33284 14356
rect 31404 14006 31432 14350
rect 33048 14272 33100 14278
rect 33048 14214 33100 14220
rect 31392 14000 31444 14006
rect 31392 13942 31444 13948
rect 31484 13932 31536 13938
rect 31484 13874 31536 13880
rect 32036 13932 32088 13938
rect 32036 13874 32088 13880
rect 31208 13796 31260 13802
rect 31208 13738 31260 13744
rect 31220 13462 31248 13738
rect 31208 13456 31260 13462
rect 31208 13398 31260 13404
rect 31496 12986 31524 13874
rect 31668 13728 31720 13734
rect 31668 13670 31720 13676
rect 31680 13258 31708 13670
rect 31944 13320 31996 13326
rect 31944 13262 31996 13268
rect 31668 13252 31720 13258
rect 31668 13194 31720 13200
rect 31484 12980 31536 12986
rect 31484 12922 31536 12928
rect 31956 12850 31984 13262
rect 31392 12844 31444 12850
rect 31392 12786 31444 12792
rect 31944 12844 31996 12850
rect 31944 12786 31996 12792
rect 31208 12776 31260 12782
rect 31208 12718 31260 12724
rect 31220 11694 31248 12718
rect 31404 12442 31432 12786
rect 31760 12708 31812 12714
rect 31760 12650 31812 12656
rect 31392 12436 31444 12442
rect 31392 12378 31444 12384
rect 31208 11688 31260 11694
rect 31208 11630 31260 11636
rect 31772 11642 31800 12650
rect 32048 12306 32076 13874
rect 32772 13864 32824 13870
rect 32772 13806 32824 13812
rect 32128 13796 32180 13802
rect 32128 13738 32180 13744
rect 32680 13796 32732 13802
rect 32680 13738 32732 13744
rect 32140 12714 32168 13738
rect 32692 13530 32720 13738
rect 32784 13530 32812 13806
rect 32680 13524 32732 13530
rect 32680 13466 32732 13472
rect 32772 13524 32824 13530
rect 32772 13466 32824 13472
rect 33060 12918 33088 14214
rect 33244 14074 33272 14350
rect 33336 14346 33364 14962
rect 34072 14618 34100 15370
rect 34348 15162 34376 15506
rect 34336 15156 34388 15162
rect 34336 15098 34388 15104
rect 34244 14952 34296 14958
rect 34244 14894 34296 14900
rect 34256 14618 34284 14894
rect 34060 14612 34112 14618
rect 34060 14554 34112 14560
rect 34244 14612 34296 14618
rect 34244 14554 34296 14560
rect 34532 14550 34560 15982
rect 34612 15972 34664 15978
rect 34612 15914 34664 15920
rect 34520 14544 34572 14550
rect 34520 14486 34572 14492
rect 34624 14414 34652 15914
rect 34796 15904 34848 15910
rect 34796 15846 34848 15852
rect 36084 15904 36136 15910
rect 36084 15846 36136 15852
rect 34808 14482 34836 15846
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 35624 15564 35676 15570
rect 35624 15506 35676 15512
rect 35636 15348 35664 15506
rect 35452 15320 35664 15348
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 35452 14618 35480 15320
rect 35594 15260 35902 15269
rect 35594 15258 35600 15260
rect 35656 15258 35680 15260
rect 35736 15258 35760 15260
rect 35816 15258 35840 15260
rect 35896 15258 35902 15260
rect 35656 15206 35658 15258
rect 35838 15206 35840 15258
rect 35594 15204 35600 15206
rect 35656 15204 35680 15206
rect 35736 15204 35760 15206
rect 35816 15204 35840 15206
rect 35896 15204 35902 15206
rect 35594 15195 35902 15204
rect 36096 15094 36124 15846
rect 36268 15360 36320 15366
rect 36268 15302 36320 15308
rect 36084 15088 36136 15094
rect 36084 15030 36136 15036
rect 36280 15026 36308 15302
rect 36268 15020 36320 15026
rect 36268 14962 36320 14968
rect 35624 14816 35676 14822
rect 35624 14758 35676 14764
rect 36176 14816 36228 14822
rect 36176 14758 36228 14764
rect 35440 14612 35492 14618
rect 35440 14554 35492 14560
rect 35636 14550 35664 14758
rect 35624 14544 35676 14550
rect 35624 14486 35676 14492
rect 34796 14476 34848 14482
rect 34796 14418 34848 14424
rect 36188 14414 36216 14758
rect 34612 14408 34664 14414
rect 34612 14350 34664 14356
rect 36176 14408 36228 14414
rect 36176 14350 36228 14356
rect 33324 14340 33376 14346
rect 33324 14282 33376 14288
rect 35594 14172 35902 14181
rect 35594 14170 35600 14172
rect 35656 14170 35680 14172
rect 35736 14170 35760 14172
rect 35816 14170 35840 14172
rect 35896 14170 35902 14172
rect 35656 14118 35658 14170
rect 35838 14118 35840 14170
rect 35594 14116 35600 14118
rect 35656 14116 35680 14118
rect 35736 14116 35760 14118
rect 35816 14116 35840 14118
rect 35896 14116 35902 14118
rect 35594 14107 35902 14116
rect 33232 14068 33284 14074
rect 33232 14010 33284 14016
rect 34796 13932 34848 13938
rect 34796 13874 34848 13880
rect 34520 13796 34572 13802
rect 34520 13738 34572 13744
rect 33784 13728 33836 13734
rect 33784 13670 33836 13676
rect 33232 13524 33284 13530
rect 33232 13466 33284 13472
rect 33244 12986 33272 13466
rect 33232 12980 33284 12986
rect 33232 12922 33284 12928
rect 33048 12912 33100 12918
rect 33048 12854 33100 12860
rect 32128 12708 32180 12714
rect 32128 12650 32180 12656
rect 33244 12434 33272 12922
rect 33796 12918 33824 13670
rect 34336 13320 34388 13326
rect 34336 13262 34388 13268
rect 34428 13320 34480 13326
rect 34428 13262 34480 13268
rect 33784 12912 33836 12918
rect 33784 12854 33836 12860
rect 33152 12406 33272 12434
rect 32036 12300 32088 12306
rect 32036 12242 32088 12248
rect 32220 12232 32272 12238
rect 32220 12174 32272 12180
rect 32036 11688 32088 11694
rect 31772 11614 31892 11642
rect 32036 11630 32088 11636
rect 31760 11552 31812 11558
rect 31760 11494 31812 11500
rect 31392 10668 31444 10674
rect 31392 10610 31444 10616
rect 31404 9178 31432 10610
rect 31772 10062 31800 11494
rect 31864 10470 31892 11614
rect 31852 10464 31904 10470
rect 31852 10406 31904 10412
rect 31864 10266 31892 10406
rect 31852 10260 31904 10266
rect 31852 10202 31904 10208
rect 31760 10056 31812 10062
rect 31760 9998 31812 10004
rect 31668 9648 31720 9654
rect 31668 9590 31720 9596
rect 31392 9172 31444 9178
rect 31392 9114 31444 9120
rect 31116 9036 31168 9042
rect 31116 8978 31168 8984
rect 31680 8634 31708 9590
rect 31760 9512 31812 9518
rect 31760 9454 31812 9460
rect 31668 8628 31720 8634
rect 31668 8570 31720 8576
rect 30840 8560 30892 8566
rect 30840 8502 30892 8508
rect 30656 7948 30708 7954
rect 30656 7890 30708 7896
rect 30288 7540 30340 7546
rect 30288 7482 30340 7488
rect 30380 7472 30432 7478
rect 30380 7414 30432 7420
rect 30288 7200 30340 7206
rect 30288 7142 30340 7148
rect 30300 6118 30328 7142
rect 30288 6112 30340 6118
rect 30288 6054 30340 6060
rect 30300 5778 30328 6054
rect 30288 5772 30340 5778
rect 30288 5714 30340 5720
rect 30392 5710 30420 7414
rect 30472 7336 30524 7342
rect 30472 7278 30524 7284
rect 30484 6458 30512 7278
rect 30852 7002 30880 8502
rect 31116 8492 31168 8498
rect 31116 8434 31168 8440
rect 31128 8090 31156 8434
rect 31116 8084 31168 8090
rect 31116 8026 31168 8032
rect 30932 8016 30984 8022
rect 31772 7970 31800 9454
rect 31852 9376 31904 9382
rect 31852 9318 31904 9324
rect 31864 8906 31892 9318
rect 32048 9042 32076 11630
rect 32232 11626 32260 12174
rect 33152 12170 33180 12406
rect 33140 12164 33192 12170
rect 33140 12106 33192 12112
rect 32772 12096 32824 12102
rect 32772 12038 32824 12044
rect 33232 12096 33284 12102
rect 33232 12038 33284 12044
rect 33968 12096 34020 12102
rect 33968 12038 34020 12044
rect 32784 11898 32812 12038
rect 33244 11898 33272 12038
rect 32772 11892 32824 11898
rect 32772 11834 32824 11840
rect 33232 11892 33284 11898
rect 33232 11834 33284 11840
rect 33048 11688 33100 11694
rect 33048 11630 33100 11636
rect 32220 11620 32272 11626
rect 32220 11562 32272 11568
rect 32404 11552 32456 11558
rect 32404 11494 32456 11500
rect 32312 11076 32364 11082
rect 32312 11018 32364 11024
rect 32324 10266 32352 11018
rect 32416 10742 32444 11494
rect 33060 11218 33088 11630
rect 33048 11212 33100 11218
rect 33048 11154 33100 11160
rect 32404 10736 32456 10742
rect 32404 10678 32456 10684
rect 33140 10736 33192 10742
rect 33140 10678 33192 10684
rect 32680 10464 32732 10470
rect 32680 10406 32732 10412
rect 32312 10260 32364 10266
rect 32312 10202 32364 10208
rect 32128 9920 32180 9926
rect 32128 9862 32180 9868
rect 32036 9036 32088 9042
rect 32036 8978 32088 8984
rect 32140 8974 32168 9862
rect 32692 9042 32720 10406
rect 33152 9994 33180 10678
rect 33244 10674 33272 11834
rect 33600 11824 33652 11830
rect 33600 11766 33652 11772
rect 33324 11688 33376 11694
rect 33324 11630 33376 11636
rect 33336 10810 33364 11630
rect 33612 11286 33640 11766
rect 33980 11354 34008 12038
rect 33968 11348 34020 11354
rect 33968 11290 34020 11296
rect 33600 11280 33652 11286
rect 33600 11222 33652 11228
rect 33612 10810 33640 11222
rect 34348 11150 34376 13262
rect 34336 11144 34388 11150
rect 34336 11086 34388 11092
rect 33692 11008 33744 11014
rect 33692 10950 33744 10956
rect 33704 10810 33732 10950
rect 33324 10804 33376 10810
rect 33324 10746 33376 10752
rect 33600 10804 33652 10810
rect 33600 10746 33652 10752
rect 33692 10804 33744 10810
rect 33692 10746 33744 10752
rect 34348 10674 34376 11086
rect 33232 10668 33284 10674
rect 33232 10610 33284 10616
rect 33692 10668 33744 10674
rect 33692 10610 33744 10616
rect 34336 10668 34388 10674
rect 34336 10610 34388 10616
rect 33600 10056 33652 10062
rect 33600 9998 33652 10004
rect 33140 9988 33192 9994
rect 33140 9930 33192 9936
rect 32956 9920 33008 9926
rect 32956 9862 33008 9868
rect 33416 9920 33468 9926
rect 33416 9862 33468 9868
rect 32968 9382 32996 9862
rect 33428 9654 33456 9862
rect 33416 9648 33468 9654
rect 33416 9590 33468 9596
rect 32956 9376 33008 9382
rect 32956 9318 33008 9324
rect 32496 9036 32548 9042
rect 32496 8978 32548 8984
rect 32680 9036 32732 9042
rect 32680 8978 32732 8984
rect 32128 8968 32180 8974
rect 32128 8910 32180 8916
rect 31852 8900 31904 8906
rect 31852 8842 31904 8848
rect 32508 8430 32536 8978
rect 32968 8974 32996 9318
rect 33612 9178 33640 9998
rect 33600 9172 33652 9178
rect 33600 9114 33652 9120
rect 33140 9036 33192 9042
rect 33140 8978 33192 8984
rect 32956 8968 33008 8974
rect 32956 8910 33008 8916
rect 32864 8492 32916 8498
rect 32864 8434 32916 8440
rect 32496 8424 32548 8430
rect 32496 8366 32548 8372
rect 32772 8424 32824 8430
rect 32772 8366 32824 8372
rect 30984 7964 31064 7970
rect 30932 7958 31064 7964
rect 30944 7942 31064 7958
rect 31772 7954 31892 7970
rect 30840 6996 30892 7002
rect 30840 6938 30892 6944
rect 31036 6866 31064 7942
rect 31760 7948 31892 7954
rect 31812 7942 31892 7948
rect 31760 7890 31812 7896
rect 31864 7342 31892 7942
rect 31852 7336 31904 7342
rect 31852 7278 31904 7284
rect 31668 6996 31720 7002
rect 31668 6938 31720 6944
rect 31680 6866 31708 6938
rect 31024 6860 31076 6866
rect 31024 6802 31076 6808
rect 31208 6860 31260 6866
rect 31208 6802 31260 6808
rect 31668 6860 31720 6866
rect 31668 6802 31720 6808
rect 30840 6656 30892 6662
rect 30840 6598 30892 6604
rect 30472 6452 30524 6458
rect 30472 6394 30524 6400
rect 30852 6322 30880 6598
rect 30840 6316 30892 6322
rect 30840 6258 30892 6264
rect 30472 6248 30524 6254
rect 30472 6190 30524 6196
rect 30380 5704 30432 5710
rect 30380 5646 30432 5652
rect 30484 5370 30512 6190
rect 31220 5778 31248 6802
rect 31300 6656 31352 6662
rect 31300 6598 31352 6604
rect 31576 6656 31628 6662
rect 31576 6598 31628 6604
rect 31312 6390 31340 6598
rect 31300 6384 31352 6390
rect 31300 6326 31352 6332
rect 31208 5772 31260 5778
rect 31208 5714 31260 5720
rect 31208 5636 31260 5642
rect 31208 5578 31260 5584
rect 30472 5364 30524 5370
rect 30472 5306 30524 5312
rect 30932 5160 30984 5166
rect 30932 5102 30984 5108
rect 30944 5030 30972 5102
rect 30932 5024 30984 5030
rect 30932 4966 30984 4972
rect 31220 4826 31248 5578
rect 31312 5234 31340 6326
rect 31588 5234 31616 6598
rect 31300 5228 31352 5234
rect 31300 5170 31352 5176
rect 31576 5228 31628 5234
rect 31576 5170 31628 5176
rect 31680 5166 31708 6802
rect 32508 5166 32536 8366
rect 32784 7750 32812 8366
rect 32772 7744 32824 7750
rect 32772 7686 32824 7692
rect 32680 7336 32732 7342
rect 32680 7278 32732 7284
rect 32692 6254 32720 7278
rect 32784 6798 32812 7686
rect 32876 6798 32904 8434
rect 33152 7954 33180 8978
rect 33600 8900 33652 8906
rect 33600 8842 33652 8848
rect 33612 8634 33640 8842
rect 33600 8628 33652 8634
rect 33600 8570 33652 8576
rect 33140 7948 33192 7954
rect 33140 7890 33192 7896
rect 32956 7812 33008 7818
rect 32956 7754 33008 7760
rect 32968 6866 32996 7754
rect 33704 7546 33732 10610
rect 34440 9738 34468 13262
rect 34532 12986 34560 13738
rect 34520 12980 34572 12986
rect 34520 12922 34572 12928
rect 34532 12374 34560 12922
rect 34520 12368 34572 12374
rect 34520 12310 34572 12316
rect 34808 12238 34836 13874
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 35594 13084 35902 13093
rect 35594 13082 35600 13084
rect 35656 13082 35680 13084
rect 35736 13082 35760 13084
rect 35816 13082 35840 13084
rect 35896 13082 35902 13084
rect 35656 13030 35658 13082
rect 35838 13030 35840 13082
rect 35594 13028 35600 13030
rect 35656 13028 35680 13030
rect 35736 13028 35760 13030
rect 35816 13028 35840 13030
rect 35896 13028 35902 13030
rect 35594 13019 35902 13028
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 34796 12232 34848 12238
rect 34796 12174 34848 12180
rect 34348 9710 34468 9738
rect 33876 9648 33928 9654
rect 33876 9590 33928 9596
rect 33888 9178 33916 9590
rect 33876 9172 33928 9178
rect 33876 9114 33928 9120
rect 33784 8968 33836 8974
rect 33784 8910 33836 8916
rect 33692 7540 33744 7546
rect 33692 7482 33744 7488
rect 33048 7336 33100 7342
rect 33048 7278 33100 7284
rect 32956 6860 33008 6866
rect 32956 6802 33008 6808
rect 32772 6792 32824 6798
rect 32772 6734 32824 6740
rect 32864 6792 32916 6798
rect 32916 6740 32996 6746
rect 32864 6734 32996 6740
rect 32876 6718 32996 6734
rect 32864 6656 32916 6662
rect 32864 6598 32916 6604
rect 32680 6248 32732 6254
rect 32680 6190 32732 6196
rect 32588 5636 32640 5642
rect 32588 5578 32640 5584
rect 31668 5160 31720 5166
rect 31668 5102 31720 5108
rect 32496 5160 32548 5166
rect 32496 5102 32548 5108
rect 32128 5024 32180 5030
rect 32128 4966 32180 4972
rect 31208 4820 31260 4826
rect 31208 4762 31260 4768
rect 31484 4752 31536 4758
rect 31484 4694 31536 4700
rect 30748 4548 30800 4554
rect 30748 4490 30800 4496
rect 30760 4146 30788 4490
rect 31496 4282 31524 4694
rect 32140 4622 32168 4966
rect 32600 4826 32628 5578
rect 32772 5568 32824 5574
rect 32772 5510 32824 5516
rect 32784 5302 32812 5510
rect 32876 5370 32904 6598
rect 32864 5364 32916 5370
rect 32864 5306 32916 5312
rect 32772 5296 32824 5302
rect 32772 5238 32824 5244
rect 32864 5160 32916 5166
rect 32864 5102 32916 5108
rect 32588 4820 32640 4826
rect 32588 4762 32640 4768
rect 32876 4690 32904 5102
rect 32864 4684 32916 4690
rect 32864 4626 32916 4632
rect 32968 4622 32996 6718
rect 33060 6662 33088 7278
rect 33508 6724 33560 6730
rect 33508 6666 33560 6672
rect 33048 6656 33100 6662
rect 33048 6598 33100 6604
rect 33520 6118 33548 6666
rect 33692 6384 33744 6390
rect 33692 6326 33744 6332
rect 33508 6112 33560 6118
rect 33508 6054 33560 6060
rect 33520 5710 33548 6054
rect 33508 5704 33560 5710
rect 33508 5646 33560 5652
rect 33704 5370 33732 6326
rect 33692 5364 33744 5370
rect 33692 5306 33744 5312
rect 33796 5234 33824 8910
rect 34348 8634 34376 9710
rect 34428 9580 34480 9586
rect 34428 9522 34480 9528
rect 34336 8628 34388 8634
rect 34336 8570 34388 8576
rect 34348 7886 34376 8570
rect 34336 7880 34388 7886
rect 34336 7822 34388 7828
rect 34152 7744 34204 7750
rect 34152 7686 34204 7692
rect 34164 6798 34192 7686
rect 34348 7546 34376 7822
rect 34336 7540 34388 7546
rect 34336 7482 34388 7488
rect 34152 6792 34204 6798
rect 34152 6734 34204 6740
rect 34244 6316 34296 6322
rect 34244 6258 34296 6264
rect 34256 5914 34284 6258
rect 34440 6118 34468 9522
rect 34808 8974 34836 12174
rect 34980 12096 35032 12102
rect 34980 12038 35032 12044
rect 34992 11830 35020 12038
rect 35594 11996 35902 12005
rect 35594 11994 35600 11996
rect 35656 11994 35680 11996
rect 35736 11994 35760 11996
rect 35816 11994 35840 11996
rect 35896 11994 35902 11996
rect 35656 11942 35658 11994
rect 35838 11942 35840 11994
rect 35594 11940 35600 11942
rect 35656 11940 35680 11942
rect 35736 11940 35760 11942
rect 35816 11940 35840 11942
rect 35896 11940 35902 11942
rect 35594 11931 35902 11940
rect 36648 11898 36676 20402
rect 36728 15904 36780 15910
rect 36728 15846 36780 15852
rect 36740 15502 36768 15846
rect 36728 15496 36780 15502
rect 36728 15438 36780 15444
rect 36832 13802 36860 22066
rect 36910 20360 36966 20369
rect 36910 20295 36912 20304
rect 36964 20295 36966 20304
rect 36912 20266 36964 20272
rect 36912 16584 36964 16590
rect 36912 16526 36964 16532
rect 36820 13796 36872 13802
rect 36820 13738 36872 13744
rect 36636 11892 36688 11898
rect 36636 11834 36688 11840
rect 34980 11824 35032 11830
rect 34980 11766 35032 11772
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 35594 10908 35902 10917
rect 35594 10906 35600 10908
rect 35656 10906 35680 10908
rect 35736 10906 35760 10908
rect 35816 10906 35840 10908
rect 35896 10906 35902 10908
rect 35656 10854 35658 10906
rect 35838 10854 35840 10906
rect 35594 10852 35600 10854
rect 35656 10852 35680 10854
rect 35736 10852 35760 10854
rect 35816 10852 35840 10854
rect 35896 10852 35902 10854
rect 35594 10843 35902 10852
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 35594 9820 35902 9829
rect 35594 9818 35600 9820
rect 35656 9818 35680 9820
rect 35736 9818 35760 9820
rect 35816 9818 35840 9820
rect 35896 9818 35902 9820
rect 35656 9766 35658 9818
rect 35838 9766 35840 9818
rect 35594 9764 35600 9766
rect 35656 9764 35680 9766
rect 35736 9764 35760 9766
rect 35816 9764 35840 9766
rect 35896 9764 35902 9766
rect 35594 9755 35902 9764
rect 36924 9518 36952 16526
rect 37016 13734 37044 27406
rect 37096 24064 37148 24070
rect 37094 24032 37096 24041
rect 37148 24032 37150 24041
rect 37094 23967 37150 23976
rect 37094 16688 37150 16697
rect 37094 16623 37150 16632
rect 37108 16454 37136 16623
rect 37096 16448 37148 16454
rect 37096 16390 37148 16396
rect 37004 13728 37056 13734
rect 37004 13670 37056 13676
rect 37096 13184 37148 13190
rect 37096 13126 37148 13132
rect 37108 13025 37136 13126
rect 37094 13016 37150 13025
rect 37094 12951 37150 12960
rect 36912 9512 36964 9518
rect 36912 9454 36964 9460
rect 36912 9376 36964 9382
rect 36910 9344 36912 9353
rect 36964 9344 36966 9353
rect 34934 9276 35242 9285
rect 36910 9279 36966 9288
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 34796 8968 34848 8974
rect 34796 8910 34848 8916
rect 34808 8498 34836 8910
rect 35594 8732 35902 8741
rect 35594 8730 35600 8732
rect 35656 8730 35680 8732
rect 35736 8730 35760 8732
rect 35816 8730 35840 8732
rect 35896 8730 35902 8732
rect 35656 8678 35658 8730
rect 35838 8678 35840 8730
rect 35594 8676 35600 8678
rect 35656 8676 35680 8678
rect 35736 8676 35760 8678
rect 35816 8676 35840 8678
rect 35896 8676 35902 8678
rect 35594 8667 35902 8676
rect 34796 8492 34848 8498
rect 34796 8434 34848 8440
rect 34612 8356 34664 8362
rect 34612 8298 34664 8304
rect 34796 8356 34848 8362
rect 34796 8298 34848 8304
rect 34624 7886 34652 8298
rect 34612 7880 34664 7886
rect 34612 7822 34664 7828
rect 34808 7478 34836 8298
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 35594 7644 35902 7653
rect 35594 7642 35600 7644
rect 35656 7642 35680 7644
rect 35736 7642 35760 7644
rect 35816 7642 35840 7644
rect 35896 7642 35902 7644
rect 35656 7590 35658 7642
rect 35838 7590 35840 7642
rect 35594 7588 35600 7590
rect 35656 7588 35680 7590
rect 35736 7588 35760 7590
rect 35816 7588 35840 7590
rect 35896 7588 35902 7590
rect 35594 7579 35902 7588
rect 34796 7472 34848 7478
rect 34796 7414 34848 7420
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 35594 6556 35902 6565
rect 35594 6554 35600 6556
rect 35656 6554 35680 6556
rect 35736 6554 35760 6556
rect 35816 6554 35840 6556
rect 35896 6554 35902 6556
rect 35656 6502 35658 6554
rect 35838 6502 35840 6554
rect 35594 6500 35600 6502
rect 35656 6500 35680 6502
rect 35736 6500 35760 6502
rect 35816 6500 35840 6502
rect 35896 6500 35902 6502
rect 35594 6491 35902 6500
rect 34428 6112 34480 6118
rect 34428 6054 34480 6060
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 34244 5908 34296 5914
rect 34244 5850 34296 5856
rect 36912 5704 36964 5710
rect 36912 5646 36964 5652
rect 37094 5672 37150 5681
rect 35594 5468 35902 5477
rect 35594 5466 35600 5468
rect 35656 5466 35680 5468
rect 35736 5466 35760 5468
rect 35816 5466 35840 5468
rect 35896 5466 35902 5468
rect 35656 5414 35658 5466
rect 35838 5414 35840 5466
rect 35594 5412 35600 5414
rect 35656 5412 35680 5414
rect 35736 5412 35760 5414
rect 35816 5412 35840 5414
rect 35896 5412 35902 5414
rect 35594 5403 35902 5412
rect 33784 5228 33836 5234
rect 33784 5170 33836 5176
rect 32128 4616 32180 4622
rect 32128 4558 32180 4564
rect 32772 4616 32824 4622
rect 32772 4558 32824 4564
rect 32956 4616 33008 4622
rect 32956 4558 33008 4564
rect 31484 4276 31536 4282
rect 31484 4218 31536 4224
rect 30748 4140 30800 4146
rect 30748 4082 30800 4088
rect 32784 3534 32812 4558
rect 33796 4078 33824 5170
rect 34796 5092 34848 5098
rect 34796 5034 34848 5040
rect 33784 4072 33836 4078
rect 33784 4014 33836 4020
rect 32772 3528 32824 3534
rect 32772 3470 32824 3476
rect 34808 2650 34836 5034
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 36924 4758 36952 5646
rect 37094 5607 37150 5616
rect 37108 5574 37136 5607
rect 37096 5568 37148 5574
rect 37096 5510 37148 5516
rect 36912 4752 36964 4758
rect 36912 4694 36964 4700
rect 35594 4380 35902 4389
rect 35594 4378 35600 4380
rect 35656 4378 35680 4380
rect 35736 4378 35760 4380
rect 35816 4378 35840 4380
rect 35896 4378 35902 4380
rect 35656 4326 35658 4378
rect 35838 4326 35840 4378
rect 35594 4324 35600 4326
rect 35656 4324 35680 4326
rect 35736 4324 35760 4326
rect 35816 4324 35840 4326
rect 35896 4324 35902 4326
rect 35594 4315 35902 4324
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 36728 3732 36780 3738
rect 36728 3674 36780 3680
rect 35594 3292 35902 3301
rect 35594 3290 35600 3292
rect 35656 3290 35680 3292
rect 35736 3290 35760 3292
rect 35816 3290 35840 3292
rect 35896 3290 35902 3292
rect 35656 3238 35658 3290
rect 35838 3238 35840 3290
rect 35594 3236 35600 3238
rect 35656 3236 35680 3238
rect 35736 3236 35760 3238
rect 35816 3236 35840 3238
rect 35896 3236 35902 3238
rect 35594 3227 35902 3236
rect 36740 3058 36768 3674
rect 36728 3052 36780 3058
rect 36728 2994 36780 3000
rect 36912 2848 36964 2854
rect 36912 2790 36964 2796
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 34796 2644 34848 2650
rect 34796 2586 34848 2592
rect 30196 2508 30248 2514
rect 30196 2450 30248 2456
rect 31760 2440 31812 2446
rect 31760 2382 31812 2388
rect 34520 2440 34572 2446
rect 34520 2382 34572 2388
rect 29000 2372 29052 2378
rect 29000 2314 29052 2320
rect 29012 800 29040 2314
rect 31772 800 31800 2382
rect 34532 800 34560 2382
rect 35594 2204 35902 2213
rect 35594 2202 35600 2204
rect 35656 2202 35680 2204
rect 35736 2202 35760 2204
rect 35816 2202 35840 2204
rect 35896 2202 35902 2204
rect 35656 2150 35658 2202
rect 35838 2150 35840 2202
rect 35594 2148 35600 2150
rect 35656 2148 35680 2150
rect 35736 2148 35760 2150
rect 35816 2148 35840 2150
rect 35896 2148 35902 2150
rect 35594 2139 35902 2148
rect 36924 2009 36952 2790
rect 37280 2304 37332 2310
rect 37280 2246 37332 2252
rect 36910 2000 36966 2009
rect 36910 1935 36966 1944
rect 37292 800 37320 2246
rect 1398 0 1454 800
rect 4158 0 4214 800
rect 6918 0 6974 800
rect 9678 0 9734 800
rect 12438 0 12494 800
rect 15198 0 15254 800
rect 17958 0 18014 800
rect 20718 0 20774 800
rect 23478 0 23534 800
rect 26238 0 26294 800
rect 28998 0 29054 800
rect 31758 0 31814 800
rect 34518 0 34574 800
rect 37278 0 37334 800
<< via2 >>
rect 1582 38664 1638 38720
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4880 38106 4936 38108
rect 4960 38106 5016 38108
rect 5040 38106 5096 38108
rect 5120 38106 5176 38108
rect 4880 38054 4926 38106
rect 4926 38054 4936 38106
rect 4960 38054 4990 38106
rect 4990 38054 5002 38106
rect 5002 38054 5016 38106
rect 5040 38054 5054 38106
rect 5054 38054 5066 38106
rect 5066 38054 5096 38106
rect 5120 38054 5130 38106
rect 5130 38054 5176 38106
rect 4880 38052 4936 38054
rect 4960 38052 5016 38054
rect 5040 38052 5096 38054
rect 5120 38052 5176 38054
rect 1582 34992 1638 35048
rect 1582 31320 1638 31376
rect 1582 27648 1638 27704
rect 1582 24012 1584 24032
rect 1584 24012 1636 24032
rect 1636 24012 1638 24032
rect 1582 23976 1638 24012
rect 1582 20324 1638 20360
rect 1582 20304 1584 20324
rect 1584 20304 1636 20324
rect 1636 20304 1638 20324
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4880 37018 4936 37020
rect 4960 37018 5016 37020
rect 5040 37018 5096 37020
rect 5120 37018 5176 37020
rect 4880 36966 4926 37018
rect 4926 36966 4936 37018
rect 4960 36966 4990 37018
rect 4990 36966 5002 37018
rect 5002 36966 5016 37018
rect 5040 36966 5054 37018
rect 5054 36966 5066 37018
rect 5066 36966 5096 37018
rect 5120 36966 5130 37018
rect 5130 36966 5176 37018
rect 4880 36964 4936 36966
rect 4960 36964 5016 36966
rect 5040 36964 5096 36966
rect 5120 36964 5176 36966
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4880 35930 4936 35932
rect 4960 35930 5016 35932
rect 5040 35930 5096 35932
rect 5120 35930 5176 35932
rect 4880 35878 4926 35930
rect 4926 35878 4936 35930
rect 4960 35878 4990 35930
rect 4990 35878 5002 35930
rect 5002 35878 5016 35930
rect 5040 35878 5054 35930
rect 5054 35878 5066 35930
rect 5066 35878 5096 35930
rect 5120 35878 5130 35930
rect 5130 35878 5176 35930
rect 4880 35876 4936 35878
rect 4960 35876 5016 35878
rect 5040 35876 5096 35878
rect 5120 35876 5176 35878
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 1582 16632 1638 16688
rect 1582 12960 1638 13016
rect 4880 34842 4936 34844
rect 4960 34842 5016 34844
rect 5040 34842 5096 34844
rect 5120 34842 5176 34844
rect 4880 34790 4926 34842
rect 4926 34790 4936 34842
rect 4960 34790 4990 34842
rect 4990 34790 5002 34842
rect 5002 34790 5016 34842
rect 5040 34790 5054 34842
rect 5054 34790 5066 34842
rect 5066 34790 5096 34842
rect 5120 34790 5130 34842
rect 5130 34790 5176 34842
rect 4880 34788 4936 34790
rect 4960 34788 5016 34790
rect 5040 34788 5096 34790
rect 5120 34788 5176 34790
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4880 33754 4936 33756
rect 4960 33754 5016 33756
rect 5040 33754 5096 33756
rect 5120 33754 5176 33756
rect 4880 33702 4926 33754
rect 4926 33702 4936 33754
rect 4960 33702 4990 33754
rect 4990 33702 5002 33754
rect 5002 33702 5016 33754
rect 5040 33702 5054 33754
rect 5054 33702 5066 33754
rect 5066 33702 5096 33754
rect 5120 33702 5130 33754
rect 5130 33702 5176 33754
rect 4880 33700 4936 33702
rect 4960 33700 5016 33702
rect 5040 33700 5096 33702
rect 5120 33700 5176 33702
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4880 32666 4936 32668
rect 4960 32666 5016 32668
rect 5040 32666 5096 32668
rect 5120 32666 5176 32668
rect 4880 32614 4926 32666
rect 4926 32614 4936 32666
rect 4960 32614 4990 32666
rect 4990 32614 5002 32666
rect 5002 32614 5016 32666
rect 5040 32614 5054 32666
rect 5054 32614 5066 32666
rect 5066 32614 5096 32666
rect 5120 32614 5130 32666
rect 5130 32614 5176 32666
rect 4880 32612 4936 32614
rect 4960 32612 5016 32614
rect 5040 32612 5096 32614
rect 5120 32612 5176 32614
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4880 31578 4936 31580
rect 4960 31578 5016 31580
rect 5040 31578 5096 31580
rect 5120 31578 5176 31580
rect 4880 31526 4926 31578
rect 4926 31526 4936 31578
rect 4960 31526 4990 31578
rect 4990 31526 5002 31578
rect 5002 31526 5016 31578
rect 5040 31526 5054 31578
rect 5054 31526 5066 31578
rect 5066 31526 5096 31578
rect 5120 31526 5130 31578
rect 5130 31526 5176 31578
rect 4880 31524 4936 31526
rect 4960 31524 5016 31526
rect 5040 31524 5096 31526
rect 5120 31524 5176 31526
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4880 30490 4936 30492
rect 4960 30490 5016 30492
rect 5040 30490 5096 30492
rect 5120 30490 5176 30492
rect 4880 30438 4926 30490
rect 4926 30438 4936 30490
rect 4960 30438 4990 30490
rect 4990 30438 5002 30490
rect 5002 30438 5016 30490
rect 5040 30438 5054 30490
rect 5054 30438 5066 30490
rect 5066 30438 5096 30490
rect 5120 30438 5130 30490
rect 5130 30438 5176 30490
rect 4880 30436 4936 30438
rect 4960 30436 5016 30438
rect 5040 30436 5096 30438
rect 5120 30436 5176 30438
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4880 29402 4936 29404
rect 4960 29402 5016 29404
rect 5040 29402 5096 29404
rect 5120 29402 5176 29404
rect 4880 29350 4926 29402
rect 4926 29350 4936 29402
rect 4960 29350 4990 29402
rect 4990 29350 5002 29402
rect 5002 29350 5016 29402
rect 5040 29350 5054 29402
rect 5054 29350 5066 29402
rect 5066 29350 5096 29402
rect 5120 29350 5130 29402
rect 5130 29350 5176 29402
rect 4880 29348 4936 29350
rect 4960 29348 5016 29350
rect 5040 29348 5096 29350
rect 5120 29348 5176 29350
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4880 28314 4936 28316
rect 4960 28314 5016 28316
rect 5040 28314 5096 28316
rect 5120 28314 5176 28316
rect 4880 28262 4926 28314
rect 4926 28262 4936 28314
rect 4960 28262 4990 28314
rect 4990 28262 5002 28314
rect 5002 28262 5016 28314
rect 5040 28262 5054 28314
rect 5054 28262 5066 28314
rect 5066 28262 5096 28314
rect 5120 28262 5130 28314
rect 5130 28262 5176 28314
rect 4880 28260 4936 28262
rect 4960 28260 5016 28262
rect 5040 28260 5096 28262
rect 5120 28260 5176 28262
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4880 27226 4936 27228
rect 4960 27226 5016 27228
rect 5040 27226 5096 27228
rect 5120 27226 5176 27228
rect 4880 27174 4926 27226
rect 4926 27174 4936 27226
rect 4960 27174 4990 27226
rect 4990 27174 5002 27226
rect 5002 27174 5016 27226
rect 5040 27174 5054 27226
rect 5054 27174 5066 27226
rect 5066 27174 5096 27226
rect 5120 27174 5130 27226
rect 5130 27174 5176 27226
rect 4880 27172 4936 27174
rect 4960 27172 5016 27174
rect 5040 27172 5096 27174
rect 5120 27172 5176 27174
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4880 26138 4936 26140
rect 4960 26138 5016 26140
rect 5040 26138 5096 26140
rect 5120 26138 5176 26140
rect 4880 26086 4926 26138
rect 4926 26086 4936 26138
rect 4960 26086 4990 26138
rect 4990 26086 5002 26138
rect 5002 26086 5016 26138
rect 5040 26086 5054 26138
rect 5054 26086 5066 26138
rect 5066 26086 5096 26138
rect 5120 26086 5130 26138
rect 5130 26086 5176 26138
rect 4880 26084 4936 26086
rect 4960 26084 5016 26086
rect 5040 26084 5096 26086
rect 5120 26084 5176 26086
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4880 25050 4936 25052
rect 4960 25050 5016 25052
rect 5040 25050 5096 25052
rect 5120 25050 5176 25052
rect 4880 24998 4926 25050
rect 4926 24998 4936 25050
rect 4960 24998 4990 25050
rect 4990 24998 5002 25050
rect 5002 24998 5016 25050
rect 5040 24998 5054 25050
rect 5054 24998 5066 25050
rect 5066 24998 5096 25050
rect 5120 24998 5130 25050
rect 5130 24998 5176 25050
rect 4880 24996 4936 24998
rect 4960 24996 5016 24998
rect 5040 24996 5096 24998
rect 5120 24996 5176 24998
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4880 23962 4936 23964
rect 4960 23962 5016 23964
rect 5040 23962 5096 23964
rect 5120 23962 5176 23964
rect 4880 23910 4926 23962
rect 4926 23910 4936 23962
rect 4960 23910 4990 23962
rect 4990 23910 5002 23962
rect 5002 23910 5016 23962
rect 5040 23910 5054 23962
rect 5054 23910 5066 23962
rect 5066 23910 5096 23962
rect 5120 23910 5130 23962
rect 5130 23910 5176 23962
rect 4880 23908 4936 23910
rect 4960 23908 5016 23910
rect 5040 23908 5096 23910
rect 5120 23908 5176 23910
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4880 22874 4936 22876
rect 4960 22874 5016 22876
rect 5040 22874 5096 22876
rect 5120 22874 5176 22876
rect 4880 22822 4926 22874
rect 4926 22822 4936 22874
rect 4960 22822 4990 22874
rect 4990 22822 5002 22874
rect 5002 22822 5016 22874
rect 5040 22822 5054 22874
rect 5054 22822 5066 22874
rect 5066 22822 5096 22874
rect 5120 22822 5130 22874
rect 5130 22822 5176 22874
rect 4880 22820 4936 22822
rect 4960 22820 5016 22822
rect 5040 22820 5096 22822
rect 5120 22820 5176 22822
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4880 21786 4936 21788
rect 4960 21786 5016 21788
rect 5040 21786 5096 21788
rect 5120 21786 5176 21788
rect 4880 21734 4926 21786
rect 4926 21734 4936 21786
rect 4960 21734 4990 21786
rect 4990 21734 5002 21786
rect 5002 21734 5016 21786
rect 5040 21734 5054 21786
rect 5054 21734 5066 21786
rect 5066 21734 5096 21786
rect 5120 21734 5130 21786
rect 5130 21734 5176 21786
rect 4880 21732 4936 21734
rect 4960 21732 5016 21734
rect 5040 21732 5096 21734
rect 5120 21732 5176 21734
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4880 20698 4936 20700
rect 4960 20698 5016 20700
rect 5040 20698 5096 20700
rect 5120 20698 5176 20700
rect 4880 20646 4926 20698
rect 4926 20646 4936 20698
rect 4960 20646 4990 20698
rect 4990 20646 5002 20698
rect 5002 20646 5016 20698
rect 5040 20646 5054 20698
rect 5054 20646 5066 20698
rect 5066 20646 5096 20698
rect 5120 20646 5130 20698
rect 5130 20646 5176 20698
rect 4880 20644 4936 20646
rect 4960 20644 5016 20646
rect 5040 20644 5096 20646
rect 5120 20644 5176 20646
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4880 19610 4936 19612
rect 4960 19610 5016 19612
rect 5040 19610 5096 19612
rect 5120 19610 5176 19612
rect 4880 19558 4926 19610
rect 4926 19558 4936 19610
rect 4960 19558 4990 19610
rect 4990 19558 5002 19610
rect 5002 19558 5016 19610
rect 5040 19558 5054 19610
rect 5054 19558 5066 19610
rect 5066 19558 5096 19610
rect 5120 19558 5130 19610
rect 5130 19558 5176 19610
rect 4880 19556 4936 19558
rect 4960 19556 5016 19558
rect 5040 19556 5096 19558
rect 5120 19556 5176 19558
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4880 18522 4936 18524
rect 4960 18522 5016 18524
rect 5040 18522 5096 18524
rect 5120 18522 5176 18524
rect 4880 18470 4926 18522
rect 4926 18470 4936 18522
rect 4960 18470 4990 18522
rect 4990 18470 5002 18522
rect 5002 18470 5016 18522
rect 5040 18470 5054 18522
rect 5054 18470 5066 18522
rect 5066 18470 5096 18522
rect 5120 18470 5130 18522
rect 5130 18470 5176 18522
rect 4880 18468 4936 18470
rect 4960 18468 5016 18470
rect 5040 18468 5096 18470
rect 5120 18468 5176 18470
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4880 17434 4936 17436
rect 4960 17434 5016 17436
rect 5040 17434 5096 17436
rect 5120 17434 5176 17436
rect 4880 17382 4926 17434
rect 4926 17382 4936 17434
rect 4960 17382 4990 17434
rect 4990 17382 5002 17434
rect 5002 17382 5016 17434
rect 5040 17382 5054 17434
rect 5054 17382 5066 17434
rect 5066 17382 5096 17434
rect 5120 17382 5130 17434
rect 5130 17382 5176 17434
rect 4880 17380 4936 17382
rect 4960 17380 5016 17382
rect 5040 17380 5096 17382
rect 5120 17380 5176 17382
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4880 16346 4936 16348
rect 4960 16346 5016 16348
rect 5040 16346 5096 16348
rect 5120 16346 5176 16348
rect 4880 16294 4926 16346
rect 4926 16294 4936 16346
rect 4960 16294 4990 16346
rect 4990 16294 5002 16346
rect 5002 16294 5016 16346
rect 5040 16294 5054 16346
rect 5054 16294 5066 16346
rect 5066 16294 5096 16346
rect 5120 16294 5130 16346
rect 5130 16294 5176 16346
rect 4880 16292 4936 16294
rect 4960 16292 5016 16294
rect 5040 16292 5096 16294
rect 5120 16292 5176 16294
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4880 15258 4936 15260
rect 4960 15258 5016 15260
rect 5040 15258 5096 15260
rect 5120 15258 5176 15260
rect 4880 15206 4926 15258
rect 4926 15206 4936 15258
rect 4960 15206 4990 15258
rect 4990 15206 5002 15258
rect 5002 15206 5016 15258
rect 5040 15206 5054 15258
rect 5054 15206 5066 15258
rect 5066 15206 5096 15258
rect 5120 15206 5130 15258
rect 5130 15206 5176 15258
rect 4880 15204 4936 15206
rect 4960 15204 5016 15206
rect 5040 15204 5096 15206
rect 5120 15204 5176 15206
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4880 14170 4936 14172
rect 4960 14170 5016 14172
rect 5040 14170 5096 14172
rect 5120 14170 5176 14172
rect 4880 14118 4926 14170
rect 4926 14118 4936 14170
rect 4960 14118 4990 14170
rect 4990 14118 5002 14170
rect 5002 14118 5016 14170
rect 5040 14118 5054 14170
rect 5054 14118 5066 14170
rect 5066 14118 5096 14170
rect 5120 14118 5130 14170
rect 5130 14118 5176 14170
rect 4880 14116 4936 14118
rect 4960 14116 5016 14118
rect 5040 14116 5096 14118
rect 5120 14116 5176 14118
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4880 13082 4936 13084
rect 4960 13082 5016 13084
rect 5040 13082 5096 13084
rect 5120 13082 5176 13084
rect 4880 13030 4926 13082
rect 4926 13030 4936 13082
rect 4960 13030 4990 13082
rect 4990 13030 5002 13082
rect 5002 13030 5016 13082
rect 5040 13030 5054 13082
rect 5054 13030 5066 13082
rect 5066 13030 5096 13082
rect 5120 13030 5130 13082
rect 5130 13030 5176 13082
rect 4880 13028 4936 13030
rect 4960 13028 5016 13030
rect 5040 13028 5096 13030
rect 5120 13028 5176 13030
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4880 11994 4936 11996
rect 4960 11994 5016 11996
rect 5040 11994 5096 11996
rect 5120 11994 5176 11996
rect 4880 11942 4926 11994
rect 4926 11942 4936 11994
rect 4960 11942 4990 11994
rect 4990 11942 5002 11994
rect 5002 11942 5016 11994
rect 5040 11942 5054 11994
rect 5054 11942 5066 11994
rect 5066 11942 5096 11994
rect 5120 11942 5130 11994
rect 5130 11942 5176 11994
rect 4880 11940 4936 11942
rect 4960 11940 5016 11942
rect 5040 11940 5096 11942
rect 5120 11940 5176 11942
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4880 10906 4936 10908
rect 4960 10906 5016 10908
rect 5040 10906 5096 10908
rect 5120 10906 5176 10908
rect 4880 10854 4926 10906
rect 4926 10854 4936 10906
rect 4960 10854 4990 10906
rect 4990 10854 5002 10906
rect 5002 10854 5016 10906
rect 5040 10854 5054 10906
rect 5054 10854 5066 10906
rect 5066 10854 5096 10906
rect 5120 10854 5130 10906
rect 5130 10854 5176 10906
rect 4880 10852 4936 10854
rect 4960 10852 5016 10854
rect 5040 10852 5096 10854
rect 5120 10852 5176 10854
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4880 9818 4936 9820
rect 4960 9818 5016 9820
rect 5040 9818 5096 9820
rect 5120 9818 5176 9820
rect 4880 9766 4926 9818
rect 4926 9766 4936 9818
rect 4960 9766 4990 9818
rect 4990 9766 5002 9818
rect 5002 9766 5016 9818
rect 5040 9766 5054 9818
rect 5054 9766 5066 9818
rect 5066 9766 5096 9818
rect 5120 9766 5130 9818
rect 5130 9766 5176 9818
rect 4880 9764 4936 9766
rect 4960 9764 5016 9766
rect 5040 9764 5096 9766
rect 5120 9764 5176 9766
rect 1582 9324 1584 9344
rect 1584 9324 1636 9344
rect 1636 9324 1638 9344
rect 1582 9288 1638 9324
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4880 8730 4936 8732
rect 4960 8730 5016 8732
rect 5040 8730 5096 8732
rect 5120 8730 5176 8732
rect 4880 8678 4926 8730
rect 4926 8678 4936 8730
rect 4960 8678 4990 8730
rect 4990 8678 5002 8730
rect 5002 8678 5016 8730
rect 5040 8678 5054 8730
rect 5054 8678 5066 8730
rect 5066 8678 5096 8730
rect 5120 8678 5130 8730
rect 5130 8678 5176 8730
rect 4880 8676 4936 8678
rect 4960 8676 5016 8678
rect 5040 8676 5096 8678
rect 5120 8676 5176 8678
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 1582 5616 1638 5672
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 15106 30252 15162 30288
rect 15106 30232 15108 30252
rect 15108 30232 15160 30252
rect 15160 30232 15162 30252
rect 12990 21936 13046 21992
rect 13266 21936 13322 21992
rect 22006 37068 22008 37088
rect 22008 37068 22060 37088
rect 22060 37068 22062 37088
rect 22006 37032 22062 37068
rect 24398 37032 24454 37088
rect 20902 30232 20958 30288
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 1582 1944 1638 2000
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 35600 38106 35656 38108
rect 35680 38106 35736 38108
rect 35760 38106 35816 38108
rect 35840 38106 35896 38108
rect 35600 38054 35646 38106
rect 35646 38054 35656 38106
rect 35680 38054 35710 38106
rect 35710 38054 35722 38106
rect 35722 38054 35736 38106
rect 35760 38054 35774 38106
rect 35774 38054 35786 38106
rect 35786 38054 35816 38106
rect 35840 38054 35850 38106
rect 35850 38054 35896 38106
rect 35600 38052 35656 38054
rect 35680 38052 35736 38054
rect 35760 38052 35816 38054
rect 35840 38052 35896 38054
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 35600 37018 35656 37020
rect 35680 37018 35736 37020
rect 35760 37018 35816 37020
rect 35840 37018 35896 37020
rect 35600 36966 35646 37018
rect 35646 36966 35656 37018
rect 35680 36966 35710 37018
rect 35710 36966 35722 37018
rect 35722 36966 35736 37018
rect 35760 36966 35774 37018
rect 35774 36966 35786 37018
rect 35786 36966 35816 37018
rect 35840 36966 35850 37018
rect 35850 36966 35896 37018
rect 35600 36964 35656 36966
rect 35680 36964 35736 36966
rect 35760 36964 35816 36966
rect 35840 36964 35896 36966
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 35600 35930 35656 35932
rect 35680 35930 35736 35932
rect 35760 35930 35816 35932
rect 35840 35930 35896 35932
rect 35600 35878 35646 35930
rect 35646 35878 35656 35930
rect 35680 35878 35710 35930
rect 35710 35878 35722 35930
rect 35722 35878 35736 35930
rect 35760 35878 35774 35930
rect 35774 35878 35786 35930
rect 35786 35878 35816 35930
rect 35840 35878 35850 35930
rect 35850 35878 35896 35930
rect 35600 35876 35656 35878
rect 35680 35876 35736 35878
rect 35760 35876 35816 35878
rect 35840 35876 35896 35878
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 35600 34842 35656 34844
rect 35680 34842 35736 34844
rect 35760 34842 35816 34844
rect 35840 34842 35896 34844
rect 35600 34790 35646 34842
rect 35646 34790 35656 34842
rect 35680 34790 35710 34842
rect 35710 34790 35722 34842
rect 35722 34790 35736 34842
rect 35760 34790 35774 34842
rect 35774 34790 35786 34842
rect 35786 34790 35816 34842
rect 35840 34790 35850 34842
rect 35850 34790 35896 34842
rect 35600 34788 35656 34790
rect 35680 34788 35736 34790
rect 35760 34788 35816 34790
rect 35840 34788 35896 34790
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 35600 33754 35656 33756
rect 35680 33754 35736 33756
rect 35760 33754 35816 33756
rect 35840 33754 35896 33756
rect 35600 33702 35646 33754
rect 35646 33702 35656 33754
rect 35680 33702 35710 33754
rect 35710 33702 35722 33754
rect 35722 33702 35736 33754
rect 35760 33702 35774 33754
rect 35774 33702 35786 33754
rect 35786 33702 35816 33754
rect 35840 33702 35850 33754
rect 35850 33702 35896 33754
rect 35600 33700 35656 33702
rect 35680 33700 35736 33702
rect 35760 33700 35816 33702
rect 35840 33700 35896 33702
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 35600 32666 35656 32668
rect 35680 32666 35736 32668
rect 35760 32666 35816 32668
rect 35840 32666 35896 32668
rect 35600 32614 35646 32666
rect 35646 32614 35656 32666
rect 35680 32614 35710 32666
rect 35710 32614 35722 32666
rect 35722 32614 35736 32666
rect 35760 32614 35774 32666
rect 35774 32614 35786 32666
rect 35786 32614 35816 32666
rect 35840 32614 35850 32666
rect 35850 32614 35896 32666
rect 35600 32612 35656 32614
rect 35680 32612 35736 32614
rect 35760 32612 35816 32614
rect 35840 32612 35896 32614
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 35600 31578 35656 31580
rect 35680 31578 35736 31580
rect 35760 31578 35816 31580
rect 35840 31578 35896 31580
rect 35600 31526 35646 31578
rect 35646 31526 35656 31578
rect 35680 31526 35710 31578
rect 35710 31526 35722 31578
rect 35722 31526 35736 31578
rect 35760 31526 35774 31578
rect 35774 31526 35786 31578
rect 35786 31526 35816 31578
rect 35840 31526 35850 31578
rect 35850 31526 35896 31578
rect 35600 31524 35656 31526
rect 35680 31524 35736 31526
rect 35760 31524 35816 31526
rect 35840 31524 35896 31526
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 35600 30490 35656 30492
rect 35680 30490 35736 30492
rect 35760 30490 35816 30492
rect 35840 30490 35896 30492
rect 35600 30438 35646 30490
rect 35646 30438 35656 30490
rect 35680 30438 35710 30490
rect 35710 30438 35722 30490
rect 35722 30438 35736 30490
rect 35760 30438 35774 30490
rect 35774 30438 35786 30490
rect 35786 30438 35816 30490
rect 35840 30438 35850 30490
rect 35850 30438 35896 30490
rect 35600 30436 35656 30438
rect 35680 30436 35736 30438
rect 35760 30436 35816 30438
rect 35840 30436 35896 30438
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 35600 29402 35656 29404
rect 35680 29402 35736 29404
rect 35760 29402 35816 29404
rect 35840 29402 35896 29404
rect 35600 29350 35646 29402
rect 35646 29350 35656 29402
rect 35680 29350 35710 29402
rect 35710 29350 35722 29402
rect 35722 29350 35736 29402
rect 35760 29350 35774 29402
rect 35774 29350 35786 29402
rect 35786 29350 35816 29402
rect 35840 29350 35850 29402
rect 35850 29350 35896 29402
rect 35600 29348 35656 29350
rect 35680 29348 35736 29350
rect 35760 29348 35816 29350
rect 35840 29348 35896 29350
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 35600 28314 35656 28316
rect 35680 28314 35736 28316
rect 35760 28314 35816 28316
rect 35840 28314 35896 28316
rect 35600 28262 35646 28314
rect 35646 28262 35656 28314
rect 35680 28262 35710 28314
rect 35710 28262 35722 28314
rect 35722 28262 35736 28314
rect 35760 28262 35774 28314
rect 35774 28262 35786 28314
rect 35786 28262 35816 28314
rect 35840 28262 35850 28314
rect 35850 28262 35896 28314
rect 35600 28260 35656 28262
rect 35680 28260 35736 28262
rect 35760 28260 35816 28262
rect 35840 28260 35896 28262
rect 35600 27226 35656 27228
rect 35680 27226 35736 27228
rect 35760 27226 35816 27228
rect 35840 27226 35896 27228
rect 35600 27174 35646 27226
rect 35646 27174 35656 27226
rect 35680 27174 35710 27226
rect 35710 27174 35722 27226
rect 35722 27174 35736 27226
rect 35760 27174 35774 27226
rect 35774 27174 35786 27226
rect 35786 27174 35816 27226
rect 35840 27174 35850 27226
rect 35850 27174 35896 27226
rect 35600 27172 35656 27174
rect 35680 27172 35736 27174
rect 35760 27172 35816 27174
rect 35840 27172 35896 27174
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 35600 26138 35656 26140
rect 35680 26138 35736 26140
rect 35760 26138 35816 26140
rect 35840 26138 35896 26140
rect 35600 26086 35646 26138
rect 35646 26086 35656 26138
rect 35680 26086 35710 26138
rect 35710 26086 35722 26138
rect 35722 26086 35736 26138
rect 35760 26086 35774 26138
rect 35774 26086 35786 26138
rect 35786 26086 35816 26138
rect 35840 26086 35850 26138
rect 35850 26086 35896 26138
rect 35600 26084 35656 26086
rect 35680 26084 35736 26086
rect 35760 26084 35816 26086
rect 35840 26084 35896 26086
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 35600 25050 35656 25052
rect 35680 25050 35736 25052
rect 35760 25050 35816 25052
rect 35840 25050 35896 25052
rect 35600 24998 35646 25050
rect 35646 24998 35656 25050
rect 35680 24998 35710 25050
rect 35710 24998 35722 25050
rect 35722 24998 35736 25050
rect 35760 24998 35774 25050
rect 35774 24998 35786 25050
rect 35786 24998 35816 25050
rect 35840 24998 35850 25050
rect 35850 24998 35896 25050
rect 35600 24996 35656 24998
rect 35680 24996 35736 24998
rect 35760 24996 35816 24998
rect 35840 24996 35896 24998
rect 35600 23962 35656 23964
rect 35680 23962 35736 23964
rect 35760 23962 35816 23964
rect 35840 23962 35896 23964
rect 35600 23910 35646 23962
rect 35646 23910 35656 23962
rect 35680 23910 35710 23962
rect 35710 23910 35722 23962
rect 35722 23910 35736 23962
rect 35760 23910 35774 23962
rect 35774 23910 35786 23962
rect 35786 23910 35816 23962
rect 35840 23910 35850 23962
rect 35850 23910 35896 23962
rect 35600 23908 35656 23910
rect 35680 23908 35736 23910
rect 35760 23908 35816 23910
rect 35840 23908 35896 23910
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 35600 22874 35656 22876
rect 35680 22874 35736 22876
rect 35760 22874 35816 22876
rect 35840 22874 35896 22876
rect 35600 22822 35646 22874
rect 35646 22822 35656 22874
rect 35680 22822 35710 22874
rect 35710 22822 35722 22874
rect 35722 22822 35736 22874
rect 35760 22822 35774 22874
rect 35774 22822 35786 22874
rect 35786 22822 35816 22874
rect 35840 22822 35850 22874
rect 35850 22822 35896 22874
rect 35600 22820 35656 22822
rect 35680 22820 35736 22822
rect 35760 22820 35816 22822
rect 35840 22820 35896 22822
rect 36910 38664 36966 38720
rect 37094 34992 37150 35048
rect 37094 31320 37150 31376
rect 37094 27648 37150 27704
rect 35600 21786 35656 21788
rect 35680 21786 35736 21788
rect 35760 21786 35816 21788
rect 35840 21786 35896 21788
rect 35600 21734 35646 21786
rect 35646 21734 35656 21786
rect 35680 21734 35710 21786
rect 35710 21734 35722 21786
rect 35722 21734 35736 21786
rect 35760 21734 35774 21786
rect 35774 21734 35786 21786
rect 35786 21734 35816 21786
rect 35840 21734 35850 21786
rect 35850 21734 35896 21786
rect 35600 21732 35656 21734
rect 35680 21732 35736 21734
rect 35760 21732 35816 21734
rect 35840 21732 35896 21734
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 35600 20698 35656 20700
rect 35680 20698 35736 20700
rect 35760 20698 35816 20700
rect 35840 20698 35896 20700
rect 35600 20646 35646 20698
rect 35646 20646 35656 20698
rect 35680 20646 35710 20698
rect 35710 20646 35722 20698
rect 35722 20646 35736 20698
rect 35760 20646 35774 20698
rect 35774 20646 35786 20698
rect 35786 20646 35816 20698
rect 35840 20646 35850 20698
rect 35850 20646 35896 20698
rect 35600 20644 35656 20646
rect 35680 20644 35736 20646
rect 35760 20644 35816 20646
rect 35840 20644 35896 20646
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 35600 19610 35656 19612
rect 35680 19610 35736 19612
rect 35760 19610 35816 19612
rect 35840 19610 35896 19612
rect 35600 19558 35646 19610
rect 35646 19558 35656 19610
rect 35680 19558 35710 19610
rect 35710 19558 35722 19610
rect 35722 19558 35736 19610
rect 35760 19558 35774 19610
rect 35774 19558 35786 19610
rect 35786 19558 35816 19610
rect 35840 19558 35850 19610
rect 35850 19558 35896 19610
rect 35600 19556 35656 19558
rect 35680 19556 35736 19558
rect 35760 19556 35816 19558
rect 35840 19556 35896 19558
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 35600 18522 35656 18524
rect 35680 18522 35736 18524
rect 35760 18522 35816 18524
rect 35840 18522 35896 18524
rect 35600 18470 35646 18522
rect 35646 18470 35656 18522
rect 35680 18470 35710 18522
rect 35710 18470 35722 18522
rect 35722 18470 35736 18522
rect 35760 18470 35774 18522
rect 35774 18470 35786 18522
rect 35786 18470 35816 18522
rect 35840 18470 35850 18522
rect 35850 18470 35896 18522
rect 35600 18468 35656 18470
rect 35680 18468 35736 18470
rect 35760 18468 35816 18470
rect 35840 18468 35896 18470
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 35600 17434 35656 17436
rect 35680 17434 35736 17436
rect 35760 17434 35816 17436
rect 35840 17434 35896 17436
rect 35600 17382 35646 17434
rect 35646 17382 35656 17434
rect 35680 17382 35710 17434
rect 35710 17382 35722 17434
rect 35722 17382 35736 17434
rect 35760 17382 35774 17434
rect 35774 17382 35786 17434
rect 35786 17382 35816 17434
rect 35840 17382 35850 17434
rect 35850 17382 35896 17434
rect 35600 17380 35656 17382
rect 35680 17380 35736 17382
rect 35760 17380 35816 17382
rect 35840 17380 35896 17382
rect 35600 16346 35656 16348
rect 35680 16346 35736 16348
rect 35760 16346 35816 16348
rect 35840 16346 35896 16348
rect 35600 16294 35646 16346
rect 35646 16294 35656 16346
rect 35680 16294 35710 16346
rect 35710 16294 35722 16346
rect 35722 16294 35736 16346
rect 35760 16294 35774 16346
rect 35774 16294 35786 16346
rect 35786 16294 35816 16346
rect 35840 16294 35850 16346
rect 35850 16294 35896 16346
rect 35600 16292 35656 16294
rect 35680 16292 35736 16294
rect 35760 16292 35816 16294
rect 35840 16292 35896 16294
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 35600 15258 35656 15260
rect 35680 15258 35736 15260
rect 35760 15258 35816 15260
rect 35840 15258 35896 15260
rect 35600 15206 35646 15258
rect 35646 15206 35656 15258
rect 35680 15206 35710 15258
rect 35710 15206 35722 15258
rect 35722 15206 35736 15258
rect 35760 15206 35774 15258
rect 35774 15206 35786 15258
rect 35786 15206 35816 15258
rect 35840 15206 35850 15258
rect 35850 15206 35896 15258
rect 35600 15204 35656 15206
rect 35680 15204 35736 15206
rect 35760 15204 35816 15206
rect 35840 15204 35896 15206
rect 35600 14170 35656 14172
rect 35680 14170 35736 14172
rect 35760 14170 35816 14172
rect 35840 14170 35896 14172
rect 35600 14118 35646 14170
rect 35646 14118 35656 14170
rect 35680 14118 35710 14170
rect 35710 14118 35722 14170
rect 35722 14118 35736 14170
rect 35760 14118 35774 14170
rect 35774 14118 35786 14170
rect 35786 14118 35816 14170
rect 35840 14118 35850 14170
rect 35850 14118 35896 14170
rect 35600 14116 35656 14118
rect 35680 14116 35736 14118
rect 35760 14116 35816 14118
rect 35840 14116 35896 14118
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 35600 13082 35656 13084
rect 35680 13082 35736 13084
rect 35760 13082 35816 13084
rect 35840 13082 35896 13084
rect 35600 13030 35646 13082
rect 35646 13030 35656 13082
rect 35680 13030 35710 13082
rect 35710 13030 35722 13082
rect 35722 13030 35736 13082
rect 35760 13030 35774 13082
rect 35774 13030 35786 13082
rect 35786 13030 35816 13082
rect 35840 13030 35850 13082
rect 35850 13030 35896 13082
rect 35600 13028 35656 13030
rect 35680 13028 35736 13030
rect 35760 13028 35816 13030
rect 35840 13028 35896 13030
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 35600 11994 35656 11996
rect 35680 11994 35736 11996
rect 35760 11994 35816 11996
rect 35840 11994 35896 11996
rect 35600 11942 35646 11994
rect 35646 11942 35656 11994
rect 35680 11942 35710 11994
rect 35710 11942 35722 11994
rect 35722 11942 35736 11994
rect 35760 11942 35774 11994
rect 35774 11942 35786 11994
rect 35786 11942 35816 11994
rect 35840 11942 35850 11994
rect 35850 11942 35896 11994
rect 35600 11940 35656 11942
rect 35680 11940 35736 11942
rect 35760 11940 35816 11942
rect 35840 11940 35896 11942
rect 36910 20324 36966 20360
rect 36910 20304 36912 20324
rect 36912 20304 36964 20324
rect 36964 20304 36966 20324
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 35600 10906 35656 10908
rect 35680 10906 35736 10908
rect 35760 10906 35816 10908
rect 35840 10906 35896 10908
rect 35600 10854 35646 10906
rect 35646 10854 35656 10906
rect 35680 10854 35710 10906
rect 35710 10854 35722 10906
rect 35722 10854 35736 10906
rect 35760 10854 35774 10906
rect 35774 10854 35786 10906
rect 35786 10854 35816 10906
rect 35840 10854 35850 10906
rect 35850 10854 35896 10906
rect 35600 10852 35656 10854
rect 35680 10852 35736 10854
rect 35760 10852 35816 10854
rect 35840 10852 35896 10854
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 35600 9818 35656 9820
rect 35680 9818 35736 9820
rect 35760 9818 35816 9820
rect 35840 9818 35896 9820
rect 35600 9766 35646 9818
rect 35646 9766 35656 9818
rect 35680 9766 35710 9818
rect 35710 9766 35722 9818
rect 35722 9766 35736 9818
rect 35760 9766 35774 9818
rect 35774 9766 35786 9818
rect 35786 9766 35816 9818
rect 35840 9766 35850 9818
rect 35850 9766 35896 9818
rect 35600 9764 35656 9766
rect 35680 9764 35736 9766
rect 35760 9764 35816 9766
rect 35840 9764 35896 9766
rect 37094 24012 37096 24032
rect 37096 24012 37148 24032
rect 37148 24012 37150 24032
rect 37094 23976 37150 24012
rect 37094 16632 37150 16688
rect 37094 12960 37150 13016
rect 36910 9324 36912 9344
rect 36912 9324 36964 9344
rect 36964 9324 36966 9344
rect 36910 9288 36966 9324
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 35600 8730 35656 8732
rect 35680 8730 35736 8732
rect 35760 8730 35816 8732
rect 35840 8730 35896 8732
rect 35600 8678 35646 8730
rect 35646 8678 35656 8730
rect 35680 8678 35710 8730
rect 35710 8678 35722 8730
rect 35722 8678 35736 8730
rect 35760 8678 35774 8730
rect 35774 8678 35786 8730
rect 35786 8678 35816 8730
rect 35840 8678 35850 8730
rect 35850 8678 35896 8730
rect 35600 8676 35656 8678
rect 35680 8676 35736 8678
rect 35760 8676 35816 8678
rect 35840 8676 35896 8678
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 35600 7642 35656 7644
rect 35680 7642 35736 7644
rect 35760 7642 35816 7644
rect 35840 7642 35896 7644
rect 35600 7590 35646 7642
rect 35646 7590 35656 7642
rect 35680 7590 35710 7642
rect 35710 7590 35722 7642
rect 35722 7590 35736 7642
rect 35760 7590 35774 7642
rect 35774 7590 35786 7642
rect 35786 7590 35816 7642
rect 35840 7590 35850 7642
rect 35850 7590 35896 7642
rect 35600 7588 35656 7590
rect 35680 7588 35736 7590
rect 35760 7588 35816 7590
rect 35840 7588 35896 7590
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 35600 6554 35656 6556
rect 35680 6554 35736 6556
rect 35760 6554 35816 6556
rect 35840 6554 35896 6556
rect 35600 6502 35646 6554
rect 35646 6502 35656 6554
rect 35680 6502 35710 6554
rect 35710 6502 35722 6554
rect 35722 6502 35736 6554
rect 35760 6502 35774 6554
rect 35774 6502 35786 6554
rect 35786 6502 35816 6554
rect 35840 6502 35850 6554
rect 35850 6502 35896 6554
rect 35600 6500 35656 6502
rect 35680 6500 35736 6502
rect 35760 6500 35816 6502
rect 35840 6500 35896 6502
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 35600 5466 35656 5468
rect 35680 5466 35736 5468
rect 35760 5466 35816 5468
rect 35840 5466 35896 5468
rect 35600 5414 35646 5466
rect 35646 5414 35656 5466
rect 35680 5414 35710 5466
rect 35710 5414 35722 5466
rect 35722 5414 35736 5466
rect 35760 5414 35774 5466
rect 35774 5414 35786 5466
rect 35786 5414 35816 5466
rect 35840 5414 35850 5466
rect 35850 5414 35896 5466
rect 35600 5412 35656 5414
rect 35680 5412 35736 5414
rect 35760 5412 35816 5414
rect 35840 5412 35896 5414
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 37094 5616 37150 5672
rect 35600 4378 35656 4380
rect 35680 4378 35736 4380
rect 35760 4378 35816 4380
rect 35840 4378 35896 4380
rect 35600 4326 35646 4378
rect 35646 4326 35656 4378
rect 35680 4326 35710 4378
rect 35710 4326 35722 4378
rect 35722 4326 35736 4378
rect 35760 4326 35774 4378
rect 35774 4326 35786 4378
rect 35786 4326 35816 4378
rect 35840 4326 35850 4378
rect 35850 4326 35896 4378
rect 35600 4324 35656 4326
rect 35680 4324 35736 4326
rect 35760 4324 35816 4326
rect 35840 4324 35896 4326
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 35600 3290 35656 3292
rect 35680 3290 35736 3292
rect 35760 3290 35816 3292
rect 35840 3290 35896 3292
rect 35600 3238 35646 3290
rect 35646 3238 35656 3290
rect 35680 3238 35710 3290
rect 35710 3238 35722 3290
rect 35722 3238 35736 3290
rect 35760 3238 35774 3290
rect 35774 3238 35786 3290
rect 35786 3238 35816 3290
rect 35840 3238 35850 3290
rect 35850 3238 35896 3290
rect 35600 3236 35656 3238
rect 35680 3236 35736 3238
rect 35760 3236 35816 3238
rect 35840 3236 35896 3238
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 35600 2202 35656 2204
rect 35680 2202 35736 2204
rect 35760 2202 35816 2204
rect 35840 2202 35896 2204
rect 35600 2150 35646 2202
rect 35646 2150 35656 2202
rect 35680 2150 35710 2202
rect 35710 2150 35722 2202
rect 35722 2150 35736 2202
rect 35760 2150 35774 2202
rect 35774 2150 35786 2202
rect 35786 2150 35816 2202
rect 35840 2150 35850 2202
rect 35850 2150 35896 2202
rect 35600 2148 35656 2150
rect 35680 2148 35736 2150
rect 35760 2148 35816 2150
rect 35840 2148 35896 2150
rect 36910 1944 36966 2000
<< metal3 >>
rect 0 38722 800 38752
rect 1577 38722 1643 38725
rect 0 38720 1643 38722
rect 0 38664 1582 38720
rect 1638 38664 1643 38720
rect 0 38662 1643 38664
rect 0 38632 800 38662
rect 1577 38659 1643 38662
rect 36905 38722 36971 38725
rect 37949 38722 38749 38752
rect 36905 38720 38749 38722
rect 36905 38664 36910 38720
rect 36966 38664 38749 38720
rect 36905 38662 38749 38664
rect 36905 38659 36971 38662
rect 4210 38656 4526 38657
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 34930 38656 35246 38657
rect 34930 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35246 38656
rect 37949 38632 38749 38662
rect 34930 38591 35246 38592
rect 4870 38112 5186 38113
rect 4870 38048 4876 38112
rect 4940 38048 4956 38112
rect 5020 38048 5036 38112
rect 5100 38048 5116 38112
rect 5180 38048 5186 38112
rect 4870 38047 5186 38048
rect 35590 38112 35906 38113
rect 35590 38048 35596 38112
rect 35660 38048 35676 38112
rect 35740 38048 35756 38112
rect 35820 38048 35836 38112
rect 35900 38048 35906 38112
rect 35590 38047 35906 38048
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 22001 37090 22067 37093
rect 24393 37090 24459 37093
rect 22001 37088 24459 37090
rect 22001 37032 22006 37088
rect 22062 37032 24398 37088
rect 24454 37032 24459 37088
rect 22001 37030 24459 37032
rect 22001 37027 22067 37030
rect 24393 37027 24459 37030
rect 4870 37024 5186 37025
rect 4870 36960 4876 37024
rect 4940 36960 4956 37024
rect 5020 36960 5036 37024
rect 5100 36960 5116 37024
rect 5180 36960 5186 37024
rect 4870 36959 5186 36960
rect 35590 37024 35906 37025
rect 35590 36960 35596 37024
rect 35660 36960 35676 37024
rect 35740 36960 35756 37024
rect 35820 36960 35836 37024
rect 35900 36960 35906 37024
rect 35590 36959 35906 36960
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 4870 35936 5186 35937
rect 4870 35872 4876 35936
rect 4940 35872 4956 35936
rect 5020 35872 5036 35936
rect 5100 35872 5116 35936
rect 5180 35872 5186 35936
rect 4870 35871 5186 35872
rect 35590 35936 35906 35937
rect 35590 35872 35596 35936
rect 35660 35872 35676 35936
rect 35740 35872 35756 35936
rect 35820 35872 35836 35936
rect 35900 35872 35906 35936
rect 35590 35871 35906 35872
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 0 35050 800 35080
rect 1577 35050 1643 35053
rect 0 35048 1643 35050
rect 0 34992 1582 35048
rect 1638 34992 1643 35048
rect 0 34990 1643 34992
rect 0 34960 800 34990
rect 1577 34987 1643 34990
rect 37089 35050 37155 35053
rect 37949 35050 38749 35080
rect 37089 35048 38749 35050
rect 37089 34992 37094 35048
rect 37150 34992 38749 35048
rect 37089 34990 38749 34992
rect 37089 34987 37155 34990
rect 37949 34960 38749 34990
rect 4870 34848 5186 34849
rect 4870 34784 4876 34848
rect 4940 34784 4956 34848
rect 5020 34784 5036 34848
rect 5100 34784 5116 34848
rect 5180 34784 5186 34848
rect 4870 34783 5186 34784
rect 35590 34848 35906 34849
rect 35590 34784 35596 34848
rect 35660 34784 35676 34848
rect 35740 34784 35756 34848
rect 35820 34784 35836 34848
rect 35900 34784 35906 34848
rect 35590 34783 35906 34784
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 4870 33760 5186 33761
rect 4870 33696 4876 33760
rect 4940 33696 4956 33760
rect 5020 33696 5036 33760
rect 5100 33696 5116 33760
rect 5180 33696 5186 33760
rect 4870 33695 5186 33696
rect 35590 33760 35906 33761
rect 35590 33696 35596 33760
rect 35660 33696 35676 33760
rect 35740 33696 35756 33760
rect 35820 33696 35836 33760
rect 35900 33696 35906 33760
rect 35590 33695 35906 33696
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 4870 32672 5186 32673
rect 4870 32608 4876 32672
rect 4940 32608 4956 32672
rect 5020 32608 5036 32672
rect 5100 32608 5116 32672
rect 5180 32608 5186 32672
rect 4870 32607 5186 32608
rect 35590 32672 35906 32673
rect 35590 32608 35596 32672
rect 35660 32608 35676 32672
rect 35740 32608 35756 32672
rect 35820 32608 35836 32672
rect 35900 32608 35906 32672
rect 35590 32607 35906 32608
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 4870 31584 5186 31585
rect 4870 31520 4876 31584
rect 4940 31520 4956 31584
rect 5020 31520 5036 31584
rect 5100 31520 5116 31584
rect 5180 31520 5186 31584
rect 4870 31519 5186 31520
rect 35590 31584 35906 31585
rect 35590 31520 35596 31584
rect 35660 31520 35676 31584
rect 35740 31520 35756 31584
rect 35820 31520 35836 31584
rect 35900 31520 35906 31584
rect 35590 31519 35906 31520
rect 0 31378 800 31408
rect 1577 31378 1643 31381
rect 0 31376 1643 31378
rect 0 31320 1582 31376
rect 1638 31320 1643 31376
rect 0 31318 1643 31320
rect 0 31288 800 31318
rect 1577 31315 1643 31318
rect 37089 31378 37155 31381
rect 37949 31378 38749 31408
rect 37089 31376 38749 31378
rect 37089 31320 37094 31376
rect 37150 31320 38749 31376
rect 37089 31318 38749 31320
rect 37089 31315 37155 31318
rect 37949 31288 38749 31318
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 4870 30496 5186 30497
rect 4870 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5186 30496
rect 4870 30431 5186 30432
rect 35590 30496 35906 30497
rect 35590 30432 35596 30496
rect 35660 30432 35676 30496
rect 35740 30432 35756 30496
rect 35820 30432 35836 30496
rect 35900 30432 35906 30496
rect 35590 30431 35906 30432
rect 15101 30290 15167 30293
rect 20897 30290 20963 30293
rect 15101 30288 20963 30290
rect 15101 30232 15106 30288
rect 15162 30232 20902 30288
rect 20958 30232 20963 30288
rect 15101 30230 20963 30232
rect 15101 30227 15167 30230
rect 20897 30227 20963 30230
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 4870 29408 5186 29409
rect 4870 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5186 29408
rect 4870 29343 5186 29344
rect 35590 29408 35906 29409
rect 35590 29344 35596 29408
rect 35660 29344 35676 29408
rect 35740 29344 35756 29408
rect 35820 29344 35836 29408
rect 35900 29344 35906 29408
rect 35590 29343 35906 29344
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 4870 28320 5186 28321
rect 4870 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5186 28320
rect 4870 28255 5186 28256
rect 35590 28320 35906 28321
rect 35590 28256 35596 28320
rect 35660 28256 35676 28320
rect 35740 28256 35756 28320
rect 35820 28256 35836 28320
rect 35900 28256 35906 28320
rect 35590 28255 35906 28256
rect 4210 27776 4526 27777
rect 0 27706 800 27736
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 1577 27706 1643 27709
rect 0 27704 1643 27706
rect 0 27648 1582 27704
rect 1638 27648 1643 27704
rect 0 27646 1643 27648
rect 0 27616 800 27646
rect 1577 27643 1643 27646
rect 37089 27706 37155 27709
rect 37949 27706 38749 27736
rect 37089 27704 38749 27706
rect 37089 27648 37094 27704
rect 37150 27648 38749 27704
rect 37089 27646 38749 27648
rect 37089 27643 37155 27646
rect 37949 27616 38749 27646
rect 4870 27232 5186 27233
rect 4870 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5186 27232
rect 4870 27167 5186 27168
rect 35590 27232 35906 27233
rect 35590 27168 35596 27232
rect 35660 27168 35676 27232
rect 35740 27168 35756 27232
rect 35820 27168 35836 27232
rect 35900 27168 35906 27232
rect 35590 27167 35906 27168
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 4870 26144 5186 26145
rect 4870 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5186 26144
rect 4870 26079 5186 26080
rect 35590 26144 35906 26145
rect 35590 26080 35596 26144
rect 35660 26080 35676 26144
rect 35740 26080 35756 26144
rect 35820 26080 35836 26144
rect 35900 26080 35906 26144
rect 35590 26079 35906 26080
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 4870 25056 5186 25057
rect 4870 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5186 25056
rect 4870 24991 5186 24992
rect 35590 25056 35906 25057
rect 35590 24992 35596 25056
rect 35660 24992 35676 25056
rect 35740 24992 35756 25056
rect 35820 24992 35836 25056
rect 35900 24992 35906 25056
rect 35590 24991 35906 24992
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 0 24034 800 24064
rect 1577 24034 1643 24037
rect 0 24032 1643 24034
rect 0 23976 1582 24032
rect 1638 23976 1643 24032
rect 0 23974 1643 23976
rect 0 23944 800 23974
rect 1577 23971 1643 23974
rect 37089 24034 37155 24037
rect 37949 24034 38749 24064
rect 37089 24032 38749 24034
rect 37089 23976 37094 24032
rect 37150 23976 38749 24032
rect 37089 23974 38749 23976
rect 37089 23971 37155 23974
rect 4870 23968 5186 23969
rect 4870 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5186 23968
rect 4870 23903 5186 23904
rect 35590 23968 35906 23969
rect 35590 23904 35596 23968
rect 35660 23904 35676 23968
rect 35740 23904 35756 23968
rect 35820 23904 35836 23968
rect 35900 23904 35906 23968
rect 37949 23944 38749 23974
rect 35590 23903 35906 23904
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 4870 22880 5186 22881
rect 4870 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5186 22880
rect 4870 22815 5186 22816
rect 35590 22880 35906 22881
rect 35590 22816 35596 22880
rect 35660 22816 35676 22880
rect 35740 22816 35756 22880
rect 35820 22816 35836 22880
rect 35900 22816 35906 22880
rect 35590 22815 35906 22816
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 12985 21994 13051 21997
rect 13261 21994 13327 21997
rect 12985 21992 13327 21994
rect 12985 21936 12990 21992
rect 13046 21936 13266 21992
rect 13322 21936 13327 21992
rect 12985 21934 13327 21936
rect 12985 21931 13051 21934
rect 13261 21931 13327 21934
rect 4870 21792 5186 21793
rect 4870 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5186 21792
rect 4870 21727 5186 21728
rect 35590 21792 35906 21793
rect 35590 21728 35596 21792
rect 35660 21728 35676 21792
rect 35740 21728 35756 21792
rect 35820 21728 35836 21792
rect 35900 21728 35906 21792
rect 35590 21727 35906 21728
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 4870 20704 5186 20705
rect 4870 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5186 20704
rect 4870 20639 5186 20640
rect 35590 20704 35906 20705
rect 35590 20640 35596 20704
rect 35660 20640 35676 20704
rect 35740 20640 35756 20704
rect 35820 20640 35836 20704
rect 35900 20640 35906 20704
rect 35590 20639 35906 20640
rect 0 20362 800 20392
rect 1577 20362 1643 20365
rect 0 20360 1643 20362
rect 0 20304 1582 20360
rect 1638 20304 1643 20360
rect 0 20302 1643 20304
rect 0 20272 800 20302
rect 1577 20299 1643 20302
rect 36905 20362 36971 20365
rect 37949 20362 38749 20392
rect 36905 20360 38749 20362
rect 36905 20304 36910 20360
rect 36966 20304 38749 20360
rect 36905 20302 38749 20304
rect 36905 20299 36971 20302
rect 37949 20272 38749 20302
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 4870 19616 5186 19617
rect 4870 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5186 19616
rect 4870 19551 5186 19552
rect 35590 19616 35906 19617
rect 35590 19552 35596 19616
rect 35660 19552 35676 19616
rect 35740 19552 35756 19616
rect 35820 19552 35836 19616
rect 35900 19552 35906 19616
rect 35590 19551 35906 19552
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 4870 18528 5186 18529
rect 4870 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5186 18528
rect 4870 18463 5186 18464
rect 35590 18528 35906 18529
rect 35590 18464 35596 18528
rect 35660 18464 35676 18528
rect 35740 18464 35756 18528
rect 35820 18464 35836 18528
rect 35900 18464 35906 18528
rect 35590 18463 35906 18464
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 4870 17440 5186 17441
rect 4870 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5186 17440
rect 4870 17375 5186 17376
rect 35590 17440 35906 17441
rect 35590 17376 35596 17440
rect 35660 17376 35676 17440
rect 35740 17376 35756 17440
rect 35820 17376 35836 17440
rect 35900 17376 35906 17440
rect 35590 17375 35906 17376
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 0 16690 800 16720
rect 1577 16690 1643 16693
rect 0 16688 1643 16690
rect 0 16632 1582 16688
rect 1638 16632 1643 16688
rect 0 16630 1643 16632
rect 0 16600 800 16630
rect 1577 16627 1643 16630
rect 37089 16690 37155 16693
rect 37949 16690 38749 16720
rect 37089 16688 38749 16690
rect 37089 16632 37094 16688
rect 37150 16632 38749 16688
rect 37089 16630 38749 16632
rect 37089 16627 37155 16630
rect 37949 16600 38749 16630
rect 4870 16352 5186 16353
rect 4870 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5186 16352
rect 4870 16287 5186 16288
rect 35590 16352 35906 16353
rect 35590 16288 35596 16352
rect 35660 16288 35676 16352
rect 35740 16288 35756 16352
rect 35820 16288 35836 16352
rect 35900 16288 35906 16352
rect 35590 16287 35906 16288
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 4870 15264 5186 15265
rect 4870 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5186 15264
rect 4870 15199 5186 15200
rect 35590 15264 35906 15265
rect 35590 15200 35596 15264
rect 35660 15200 35676 15264
rect 35740 15200 35756 15264
rect 35820 15200 35836 15264
rect 35900 15200 35906 15264
rect 35590 15199 35906 15200
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 4870 14176 5186 14177
rect 4870 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5186 14176
rect 4870 14111 5186 14112
rect 35590 14176 35906 14177
rect 35590 14112 35596 14176
rect 35660 14112 35676 14176
rect 35740 14112 35756 14176
rect 35820 14112 35836 14176
rect 35900 14112 35906 14176
rect 35590 14111 35906 14112
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 4870 13088 5186 13089
rect 0 13018 800 13048
rect 4870 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5186 13088
rect 4870 13023 5186 13024
rect 35590 13088 35906 13089
rect 35590 13024 35596 13088
rect 35660 13024 35676 13088
rect 35740 13024 35756 13088
rect 35820 13024 35836 13088
rect 35900 13024 35906 13088
rect 35590 13023 35906 13024
rect 1577 13018 1643 13021
rect 0 13016 1643 13018
rect 0 12960 1582 13016
rect 1638 12960 1643 13016
rect 0 12958 1643 12960
rect 0 12928 800 12958
rect 1577 12955 1643 12958
rect 37089 13018 37155 13021
rect 37949 13018 38749 13048
rect 37089 13016 38749 13018
rect 37089 12960 37094 13016
rect 37150 12960 38749 13016
rect 37089 12958 38749 12960
rect 37089 12955 37155 12958
rect 37949 12928 38749 12958
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 4870 12000 5186 12001
rect 4870 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5186 12000
rect 4870 11935 5186 11936
rect 35590 12000 35906 12001
rect 35590 11936 35596 12000
rect 35660 11936 35676 12000
rect 35740 11936 35756 12000
rect 35820 11936 35836 12000
rect 35900 11936 35906 12000
rect 35590 11935 35906 11936
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 4870 10912 5186 10913
rect 4870 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5186 10912
rect 4870 10847 5186 10848
rect 35590 10912 35906 10913
rect 35590 10848 35596 10912
rect 35660 10848 35676 10912
rect 35740 10848 35756 10912
rect 35820 10848 35836 10912
rect 35900 10848 35906 10912
rect 35590 10847 35906 10848
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 4870 9824 5186 9825
rect 4870 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5186 9824
rect 4870 9759 5186 9760
rect 35590 9824 35906 9825
rect 35590 9760 35596 9824
rect 35660 9760 35676 9824
rect 35740 9760 35756 9824
rect 35820 9760 35836 9824
rect 35900 9760 35906 9824
rect 35590 9759 35906 9760
rect 0 9346 800 9376
rect 1577 9346 1643 9349
rect 0 9344 1643 9346
rect 0 9288 1582 9344
rect 1638 9288 1643 9344
rect 0 9286 1643 9288
rect 0 9256 800 9286
rect 1577 9283 1643 9286
rect 36905 9346 36971 9349
rect 37949 9346 38749 9376
rect 36905 9344 38749 9346
rect 36905 9288 36910 9344
rect 36966 9288 38749 9344
rect 36905 9286 38749 9288
rect 36905 9283 36971 9286
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 37949 9256 38749 9286
rect 34930 9215 35246 9216
rect 4870 8736 5186 8737
rect 4870 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5186 8736
rect 4870 8671 5186 8672
rect 35590 8736 35906 8737
rect 35590 8672 35596 8736
rect 35660 8672 35676 8736
rect 35740 8672 35756 8736
rect 35820 8672 35836 8736
rect 35900 8672 35906 8736
rect 35590 8671 35906 8672
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 4870 7648 5186 7649
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 4870 7583 5186 7584
rect 35590 7648 35906 7649
rect 35590 7584 35596 7648
rect 35660 7584 35676 7648
rect 35740 7584 35756 7648
rect 35820 7584 35836 7648
rect 35900 7584 35906 7648
rect 35590 7583 35906 7584
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 35590 6560 35906 6561
rect 35590 6496 35596 6560
rect 35660 6496 35676 6560
rect 35740 6496 35756 6560
rect 35820 6496 35836 6560
rect 35900 6496 35906 6560
rect 35590 6495 35906 6496
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 0 5674 800 5704
rect 1577 5674 1643 5677
rect 0 5672 1643 5674
rect 0 5616 1582 5672
rect 1638 5616 1643 5672
rect 0 5614 1643 5616
rect 0 5584 800 5614
rect 1577 5611 1643 5614
rect 37089 5674 37155 5677
rect 37949 5674 38749 5704
rect 37089 5672 38749 5674
rect 37089 5616 37094 5672
rect 37150 5616 38749 5672
rect 37089 5614 38749 5616
rect 37089 5611 37155 5614
rect 37949 5584 38749 5614
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 4870 5407 5186 5408
rect 35590 5472 35906 5473
rect 35590 5408 35596 5472
rect 35660 5408 35676 5472
rect 35740 5408 35756 5472
rect 35820 5408 35836 5472
rect 35900 5408 35906 5472
rect 35590 5407 35906 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 4870 4319 5186 4320
rect 35590 4384 35906 4385
rect 35590 4320 35596 4384
rect 35660 4320 35676 4384
rect 35740 4320 35756 4384
rect 35820 4320 35836 4384
rect 35900 4320 35906 4384
rect 35590 4319 35906 4320
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 35590 3296 35906 3297
rect 35590 3232 35596 3296
rect 35660 3232 35676 3296
rect 35740 3232 35756 3296
rect 35820 3232 35836 3296
rect 35900 3232 35906 3296
rect 35590 3231 35906 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 4870 2208 5186 2209
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 4870 2143 5186 2144
rect 35590 2208 35906 2209
rect 35590 2144 35596 2208
rect 35660 2144 35676 2208
rect 35740 2144 35756 2208
rect 35820 2144 35836 2208
rect 35900 2144 35906 2208
rect 35590 2143 35906 2144
rect 0 2002 800 2032
rect 1577 2002 1643 2005
rect 0 2000 1643 2002
rect 0 1944 1582 2000
rect 1638 1944 1643 2000
rect 0 1942 1643 1944
rect 0 1912 800 1942
rect 1577 1939 1643 1942
rect 36905 2002 36971 2005
rect 37949 2002 38749 2032
rect 36905 2000 38749 2002
rect 36905 1944 36910 2000
rect 36966 1944 38749 2000
rect 36905 1942 38749 1944
rect 36905 1939 36971 1942
rect 37949 1912 38749 1942
<< via3 >>
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 4876 38108 4940 38112
rect 4876 38052 4880 38108
rect 4880 38052 4936 38108
rect 4936 38052 4940 38108
rect 4876 38048 4940 38052
rect 4956 38108 5020 38112
rect 4956 38052 4960 38108
rect 4960 38052 5016 38108
rect 5016 38052 5020 38108
rect 4956 38048 5020 38052
rect 5036 38108 5100 38112
rect 5036 38052 5040 38108
rect 5040 38052 5096 38108
rect 5096 38052 5100 38108
rect 5036 38048 5100 38052
rect 5116 38108 5180 38112
rect 5116 38052 5120 38108
rect 5120 38052 5176 38108
rect 5176 38052 5180 38108
rect 5116 38048 5180 38052
rect 35596 38108 35660 38112
rect 35596 38052 35600 38108
rect 35600 38052 35656 38108
rect 35656 38052 35660 38108
rect 35596 38048 35660 38052
rect 35676 38108 35740 38112
rect 35676 38052 35680 38108
rect 35680 38052 35736 38108
rect 35736 38052 35740 38108
rect 35676 38048 35740 38052
rect 35756 38108 35820 38112
rect 35756 38052 35760 38108
rect 35760 38052 35816 38108
rect 35816 38052 35820 38108
rect 35756 38048 35820 38052
rect 35836 38108 35900 38112
rect 35836 38052 35840 38108
rect 35840 38052 35896 38108
rect 35896 38052 35900 38108
rect 35836 38048 35900 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 4876 37020 4940 37024
rect 4876 36964 4880 37020
rect 4880 36964 4936 37020
rect 4936 36964 4940 37020
rect 4876 36960 4940 36964
rect 4956 37020 5020 37024
rect 4956 36964 4960 37020
rect 4960 36964 5016 37020
rect 5016 36964 5020 37020
rect 4956 36960 5020 36964
rect 5036 37020 5100 37024
rect 5036 36964 5040 37020
rect 5040 36964 5096 37020
rect 5096 36964 5100 37020
rect 5036 36960 5100 36964
rect 5116 37020 5180 37024
rect 5116 36964 5120 37020
rect 5120 36964 5176 37020
rect 5176 36964 5180 37020
rect 5116 36960 5180 36964
rect 35596 37020 35660 37024
rect 35596 36964 35600 37020
rect 35600 36964 35656 37020
rect 35656 36964 35660 37020
rect 35596 36960 35660 36964
rect 35676 37020 35740 37024
rect 35676 36964 35680 37020
rect 35680 36964 35736 37020
rect 35736 36964 35740 37020
rect 35676 36960 35740 36964
rect 35756 37020 35820 37024
rect 35756 36964 35760 37020
rect 35760 36964 35816 37020
rect 35816 36964 35820 37020
rect 35756 36960 35820 36964
rect 35836 37020 35900 37024
rect 35836 36964 35840 37020
rect 35840 36964 35896 37020
rect 35896 36964 35900 37020
rect 35836 36960 35900 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 4876 35932 4940 35936
rect 4876 35876 4880 35932
rect 4880 35876 4936 35932
rect 4936 35876 4940 35932
rect 4876 35872 4940 35876
rect 4956 35932 5020 35936
rect 4956 35876 4960 35932
rect 4960 35876 5016 35932
rect 5016 35876 5020 35932
rect 4956 35872 5020 35876
rect 5036 35932 5100 35936
rect 5036 35876 5040 35932
rect 5040 35876 5096 35932
rect 5096 35876 5100 35932
rect 5036 35872 5100 35876
rect 5116 35932 5180 35936
rect 5116 35876 5120 35932
rect 5120 35876 5176 35932
rect 5176 35876 5180 35932
rect 5116 35872 5180 35876
rect 35596 35932 35660 35936
rect 35596 35876 35600 35932
rect 35600 35876 35656 35932
rect 35656 35876 35660 35932
rect 35596 35872 35660 35876
rect 35676 35932 35740 35936
rect 35676 35876 35680 35932
rect 35680 35876 35736 35932
rect 35736 35876 35740 35932
rect 35676 35872 35740 35876
rect 35756 35932 35820 35936
rect 35756 35876 35760 35932
rect 35760 35876 35816 35932
rect 35816 35876 35820 35932
rect 35756 35872 35820 35876
rect 35836 35932 35900 35936
rect 35836 35876 35840 35932
rect 35840 35876 35896 35932
rect 35896 35876 35900 35932
rect 35836 35872 35900 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 4876 34844 4940 34848
rect 4876 34788 4880 34844
rect 4880 34788 4936 34844
rect 4936 34788 4940 34844
rect 4876 34784 4940 34788
rect 4956 34844 5020 34848
rect 4956 34788 4960 34844
rect 4960 34788 5016 34844
rect 5016 34788 5020 34844
rect 4956 34784 5020 34788
rect 5036 34844 5100 34848
rect 5036 34788 5040 34844
rect 5040 34788 5096 34844
rect 5096 34788 5100 34844
rect 5036 34784 5100 34788
rect 5116 34844 5180 34848
rect 5116 34788 5120 34844
rect 5120 34788 5176 34844
rect 5176 34788 5180 34844
rect 5116 34784 5180 34788
rect 35596 34844 35660 34848
rect 35596 34788 35600 34844
rect 35600 34788 35656 34844
rect 35656 34788 35660 34844
rect 35596 34784 35660 34788
rect 35676 34844 35740 34848
rect 35676 34788 35680 34844
rect 35680 34788 35736 34844
rect 35736 34788 35740 34844
rect 35676 34784 35740 34788
rect 35756 34844 35820 34848
rect 35756 34788 35760 34844
rect 35760 34788 35816 34844
rect 35816 34788 35820 34844
rect 35756 34784 35820 34788
rect 35836 34844 35900 34848
rect 35836 34788 35840 34844
rect 35840 34788 35896 34844
rect 35896 34788 35900 34844
rect 35836 34784 35900 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 4876 33756 4940 33760
rect 4876 33700 4880 33756
rect 4880 33700 4936 33756
rect 4936 33700 4940 33756
rect 4876 33696 4940 33700
rect 4956 33756 5020 33760
rect 4956 33700 4960 33756
rect 4960 33700 5016 33756
rect 5016 33700 5020 33756
rect 4956 33696 5020 33700
rect 5036 33756 5100 33760
rect 5036 33700 5040 33756
rect 5040 33700 5096 33756
rect 5096 33700 5100 33756
rect 5036 33696 5100 33700
rect 5116 33756 5180 33760
rect 5116 33700 5120 33756
rect 5120 33700 5176 33756
rect 5176 33700 5180 33756
rect 5116 33696 5180 33700
rect 35596 33756 35660 33760
rect 35596 33700 35600 33756
rect 35600 33700 35656 33756
rect 35656 33700 35660 33756
rect 35596 33696 35660 33700
rect 35676 33756 35740 33760
rect 35676 33700 35680 33756
rect 35680 33700 35736 33756
rect 35736 33700 35740 33756
rect 35676 33696 35740 33700
rect 35756 33756 35820 33760
rect 35756 33700 35760 33756
rect 35760 33700 35816 33756
rect 35816 33700 35820 33756
rect 35756 33696 35820 33700
rect 35836 33756 35900 33760
rect 35836 33700 35840 33756
rect 35840 33700 35896 33756
rect 35896 33700 35900 33756
rect 35836 33696 35900 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 4876 32668 4940 32672
rect 4876 32612 4880 32668
rect 4880 32612 4936 32668
rect 4936 32612 4940 32668
rect 4876 32608 4940 32612
rect 4956 32668 5020 32672
rect 4956 32612 4960 32668
rect 4960 32612 5016 32668
rect 5016 32612 5020 32668
rect 4956 32608 5020 32612
rect 5036 32668 5100 32672
rect 5036 32612 5040 32668
rect 5040 32612 5096 32668
rect 5096 32612 5100 32668
rect 5036 32608 5100 32612
rect 5116 32668 5180 32672
rect 5116 32612 5120 32668
rect 5120 32612 5176 32668
rect 5176 32612 5180 32668
rect 5116 32608 5180 32612
rect 35596 32668 35660 32672
rect 35596 32612 35600 32668
rect 35600 32612 35656 32668
rect 35656 32612 35660 32668
rect 35596 32608 35660 32612
rect 35676 32668 35740 32672
rect 35676 32612 35680 32668
rect 35680 32612 35736 32668
rect 35736 32612 35740 32668
rect 35676 32608 35740 32612
rect 35756 32668 35820 32672
rect 35756 32612 35760 32668
rect 35760 32612 35816 32668
rect 35816 32612 35820 32668
rect 35756 32608 35820 32612
rect 35836 32668 35900 32672
rect 35836 32612 35840 32668
rect 35840 32612 35896 32668
rect 35896 32612 35900 32668
rect 35836 32608 35900 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 4876 31580 4940 31584
rect 4876 31524 4880 31580
rect 4880 31524 4936 31580
rect 4936 31524 4940 31580
rect 4876 31520 4940 31524
rect 4956 31580 5020 31584
rect 4956 31524 4960 31580
rect 4960 31524 5016 31580
rect 5016 31524 5020 31580
rect 4956 31520 5020 31524
rect 5036 31580 5100 31584
rect 5036 31524 5040 31580
rect 5040 31524 5096 31580
rect 5096 31524 5100 31580
rect 5036 31520 5100 31524
rect 5116 31580 5180 31584
rect 5116 31524 5120 31580
rect 5120 31524 5176 31580
rect 5176 31524 5180 31580
rect 5116 31520 5180 31524
rect 35596 31580 35660 31584
rect 35596 31524 35600 31580
rect 35600 31524 35656 31580
rect 35656 31524 35660 31580
rect 35596 31520 35660 31524
rect 35676 31580 35740 31584
rect 35676 31524 35680 31580
rect 35680 31524 35736 31580
rect 35736 31524 35740 31580
rect 35676 31520 35740 31524
rect 35756 31580 35820 31584
rect 35756 31524 35760 31580
rect 35760 31524 35816 31580
rect 35816 31524 35820 31580
rect 35756 31520 35820 31524
rect 35836 31580 35900 31584
rect 35836 31524 35840 31580
rect 35840 31524 35896 31580
rect 35896 31524 35900 31580
rect 35836 31520 35900 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 4876 30492 4940 30496
rect 4876 30436 4880 30492
rect 4880 30436 4936 30492
rect 4936 30436 4940 30492
rect 4876 30432 4940 30436
rect 4956 30492 5020 30496
rect 4956 30436 4960 30492
rect 4960 30436 5016 30492
rect 5016 30436 5020 30492
rect 4956 30432 5020 30436
rect 5036 30492 5100 30496
rect 5036 30436 5040 30492
rect 5040 30436 5096 30492
rect 5096 30436 5100 30492
rect 5036 30432 5100 30436
rect 5116 30492 5180 30496
rect 5116 30436 5120 30492
rect 5120 30436 5176 30492
rect 5176 30436 5180 30492
rect 5116 30432 5180 30436
rect 35596 30492 35660 30496
rect 35596 30436 35600 30492
rect 35600 30436 35656 30492
rect 35656 30436 35660 30492
rect 35596 30432 35660 30436
rect 35676 30492 35740 30496
rect 35676 30436 35680 30492
rect 35680 30436 35736 30492
rect 35736 30436 35740 30492
rect 35676 30432 35740 30436
rect 35756 30492 35820 30496
rect 35756 30436 35760 30492
rect 35760 30436 35816 30492
rect 35816 30436 35820 30492
rect 35756 30432 35820 30436
rect 35836 30492 35900 30496
rect 35836 30436 35840 30492
rect 35840 30436 35896 30492
rect 35896 30436 35900 30492
rect 35836 30432 35900 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 4876 29404 4940 29408
rect 4876 29348 4880 29404
rect 4880 29348 4936 29404
rect 4936 29348 4940 29404
rect 4876 29344 4940 29348
rect 4956 29404 5020 29408
rect 4956 29348 4960 29404
rect 4960 29348 5016 29404
rect 5016 29348 5020 29404
rect 4956 29344 5020 29348
rect 5036 29404 5100 29408
rect 5036 29348 5040 29404
rect 5040 29348 5096 29404
rect 5096 29348 5100 29404
rect 5036 29344 5100 29348
rect 5116 29404 5180 29408
rect 5116 29348 5120 29404
rect 5120 29348 5176 29404
rect 5176 29348 5180 29404
rect 5116 29344 5180 29348
rect 35596 29404 35660 29408
rect 35596 29348 35600 29404
rect 35600 29348 35656 29404
rect 35656 29348 35660 29404
rect 35596 29344 35660 29348
rect 35676 29404 35740 29408
rect 35676 29348 35680 29404
rect 35680 29348 35736 29404
rect 35736 29348 35740 29404
rect 35676 29344 35740 29348
rect 35756 29404 35820 29408
rect 35756 29348 35760 29404
rect 35760 29348 35816 29404
rect 35816 29348 35820 29404
rect 35756 29344 35820 29348
rect 35836 29404 35900 29408
rect 35836 29348 35840 29404
rect 35840 29348 35896 29404
rect 35896 29348 35900 29404
rect 35836 29344 35900 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 4876 28316 4940 28320
rect 4876 28260 4880 28316
rect 4880 28260 4936 28316
rect 4936 28260 4940 28316
rect 4876 28256 4940 28260
rect 4956 28316 5020 28320
rect 4956 28260 4960 28316
rect 4960 28260 5016 28316
rect 5016 28260 5020 28316
rect 4956 28256 5020 28260
rect 5036 28316 5100 28320
rect 5036 28260 5040 28316
rect 5040 28260 5096 28316
rect 5096 28260 5100 28316
rect 5036 28256 5100 28260
rect 5116 28316 5180 28320
rect 5116 28260 5120 28316
rect 5120 28260 5176 28316
rect 5176 28260 5180 28316
rect 5116 28256 5180 28260
rect 35596 28316 35660 28320
rect 35596 28260 35600 28316
rect 35600 28260 35656 28316
rect 35656 28260 35660 28316
rect 35596 28256 35660 28260
rect 35676 28316 35740 28320
rect 35676 28260 35680 28316
rect 35680 28260 35736 28316
rect 35736 28260 35740 28316
rect 35676 28256 35740 28260
rect 35756 28316 35820 28320
rect 35756 28260 35760 28316
rect 35760 28260 35816 28316
rect 35816 28260 35820 28316
rect 35756 28256 35820 28260
rect 35836 28316 35900 28320
rect 35836 28260 35840 28316
rect 35840 28260 35896 28316
rect 35896 28260 35900 28316
rect 35836 28256 35900 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 4876 27228 4940 27232
rect 4876 27172 4880 27228
rect 4880 27172 4936 27228
rect 4936 27172 4940 27228
rect 4876 27168 4940 27172
rect 4956 27228 5020 27232
rect 4956 27172 4960 27228
rect 4960 27172 5016 27228
rect 5016 27172 5020 27228
rect 4956 27168 5020 27172
rect 5036 27228 5100 27232
rect 5036 27172 5040 27228
rect 5040 27172 5096 27228
rect 5096 27172 5100 27228
rect 5036 27168 5100 27172
rect 5116 27228 5180 27232
rect 5116 27172 5120 27228
rect 5120 27172 5176 27228
rect 5176 27172 5180 27228
rect 5116 27168 5180 27172
rect 35596 27228 35660 27232
rect 35596 27172 35600 27228
rect 35600 27172 35656 27228
rect 35656 27172 35660 27228
rect 35596 27168 35660 27172
rect 35676 27228 35740 27232
rect 35676 27172 35680 27228
rect 35680 27172 35736 27228
rect 35736 27172 35740 27228
rect 35676 27168 35740 27172
rect 35756 27228 35820 27232
rect 35756 27172 35760 27228
rect 35760 27172 35816 27228
rect 35816 27172 35820 27228
rect 35756 27168 35820 27172
rect 35836 27228 35900 27232
rect 35836 27172 35840 27228
rect 35840 27172 35896 27228
rect 35896 27172 35900 27228
rect 35836 27168 35900 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 4876 26140 4940 26144
rect 4876 26084 4880 26140
rect 4880 26084 4936 26140
rect 4936 26084 4940 26140
rect 4876 26080 4940 26084
rect 4956 26140 5020 26144
rect 4956 26084 4960 26140
rect 4960 26084 5016 26140
rect 5016 26084 5020 26140
rect 4956 26080 5020 26084
rect 5036 26140 5100 26144
rect 5036 26084 5040 26140
rect 5040 26084 5096 26140
rect 5096 26084 5100 26140
rect 5036 26080 5100 26084
rect 5116 26140 5180 26144
rect 5116 26084 5120 26140
rect 5120 26084 5176 26140
rect 5176 26084 5180 26140
rect 5116 26080 5180 26084
rect 35596 26140 35660 26144
rect 35596 26084 35600 26140
rect 35600 26084 35656 26140
rect 35656 26084 35660 26140
rect 35596 26080 35660 26084
rect 35676 26140 35740 26144
rect 35676 26084 35680 26140
rect 35680 26084 35736 26140
rect 35736 26084 35740 26140
rect 35676 26080 35740 26084
rect 35756 26140 35820 26144
rect 35756 26084 35760 26140
rect 35760 26084 35816 26140
rect 35816 26084 35820 26140
rect 35756 26080 35820 26084
rect 35836 26140 35900 26144
rect 35836 26084 35840 26140
rect 35840 26084 35896 26140
rect 35896 26084 35900 26140
rect 35836 26080 35900 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 4876 25052 4940 25056
rect 4876 24996 4880 25052
rect 4880 24996 4936 25052
rect 4936 24996 4940 25052
rect 4876 24992 4940 24996
rect 4956 25052 5020 25056
rect 4956 24996 4960 25052
rect 4960 24996 5016 25052
rect 5016 24996 5020 25052
rect 4956 24992 5020 24996
rect 5036 25052 5100 25056
rect 5036 24996 5040 25052
rect 5040 24996 5096 25052
rect 5096 24996 5100 25052
rect 5036 24992 5100 24996
rect 5116 25052 5180 25056
rect 5116 24996 5120 25052
rect 5120 24996 5176 25052
rect 5176 24996 5180 25052
rect 5116 24992 5180 24996
rect 35596 25052 35660 25056
rect 35596 24996 35600 25052
rect 35600 24996 35656 25052
rect 35656 24996 35660 25052
rect 35596 24992 35660 24996
rect 35676 25052 35740 25056
rect 35676 24996 35680 25052
rect 35680 24996 35736 25052
rect 35736 24996 35740 25052
rect 35676 24992 35740 24996
rect 35756 25052 35820 25056
rect 35756 24996 35760 25052
rect 35760 24996 35816 25052
rect 35816 24996 35820 25052
rect 35756 24992 35820 24996
rect 35836 25052 35900 25056
rect 35836 24996 35840 25052
rect 35840 24996 35896 25052
rect 35896 24996 35900 25052
rect 35836 24992 35900 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 4876 23964 4940 23968
rect 4876 23908 4880 23964
rect 4880 23908 4936 23964
rect 4936 23908 4940 23964
rect 4876 23904 4940 23908
rect 4956 23964 5020 23968
rect 4956 23908 4960 23964
rect 4960 23908 5016 23964
rect 5016 23908 5020 23964
rect 4956 23904 5020 23908
rect 5036 23964 5100 23968
rect 5036 23908 5040 23964
rect 5040 23908 5096 23964
rect 5096 23908 5100 23964
rect 5036 23904 5100 23908
rect 5116 23964 5180 23968
rect 5116 23908 5120 23964
rect 5120 23908 5176 23964
rect 5176 23908 5180 23964
rect 5116 23904 5180 23908
rect 35596 23964 35660 23968
rect 35596 23908 35600 23964
rect 35600 23908 35656 23964
rect 35656 23908 35660 23964
rect 35596 23904 35660 23908
rect 35676 23964 35740 23968
rect 35676 23908 35680 23964
rect 35680 23908 35736 23964
rect 35736 23908 35740 23964
rect 35676 23904 35740 23908
rect 35756 23964 35820 23968
rect 35756 23908 35760 23964
rect 35760 23908 35816 23964
rect 35816 23908 35820 23964
rect 35756 23904 35820 23908
rect 35836 23964 35900 23968
rect 35836 23908 35840 23964
rect 35840 23908 35896 23964
rect 35896 23908 35900 23964
rect 35836 23904 35900 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 4876 22876 4940 22880
rect 4876 22820 4880 22876
rect 4880 22820 4936 22876
rect 4936 22820 4940 22876
rect 4876 22816 4940 22820
rect 4956 22876 5020 22880
rect 4956 22820 4960 22876
rect 4960 22820 5016 22876
rect 5016 22820 5020 22876
rect 4956 22816 5020 22820
rect 5036 22876 5100 22880
rect 5036 22820 5040 22876
rect 5040 22820 5096 22876
rect 5096 22820 5100 22876
rect 5036 22816 5100 22820
rect 5116 22876 5180 22880
rect 5116 22820 5120 22876
rect 5120 22820 5176 22876
rect 5176 22820 5180 22876
rect 5116 22816 5180 22820
rect 35596 22876 35660 22880
rect 35596 22820 35600 22876
rect 35600 22820 35656 22876
rect 35656 22820 35660 22876
rect 35596 22816 35660 22820
rect 35676 22876 35740 22880
rect 35676 22820 35680 22876
rect 35680 22820 35736 22876
rect 35736 22820 35740 22876
rect 35676 22816 35740 22820
rect 35756 22876 35820 22880
rect 35756 22820 35760 22876
rect 35760 22820 35816 22876
rect 35816 22820 35820 22876
rect 35756 22816 35820 22820
rect 35836 22876 35900 22880
rect 35836 22820 35840 22876
rect 35840 22820 35896 22876
rect 35896 22820 35900 22876
rect 35836 22816 35900 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 4876 21788 4940 21792
rect 4876 21732 4880 21788
rect 4880 21732 4936 21788
rect 4936 21732 4940 21788
rect 4876 21728 4940 21732
rect 4956 21788 5020 21792
rect 4956 21732 4960 21788
rect 4960 21732 5016 21788
rect 5016 21732 5020 21788
rect 4956 21728 5020 21732
rect 5036 21788 5100 21792
rect 5036 21732 5040 21788
rect 5040 21732 5096 21788
rect 5096 21732 5100 21788
rect 5036 21728 5100 21732
rect 5116 21788 5180 21792
rect 5116 21732 5120 21788
rect 5120 21732 5176 21788
rect 5176 21732 5180 21788
rect 5116 21728 5180 21732
rect 35596 21788 35660 21792
rect 35596 21732 35600 21788
rect 35600 21732 35656 21788
rect 35656 21732 35660 21788
rect 35596 21728 35660 21732
rect 35676 21788 35740 21792
rect 35676 21732 35680 21788
rect 35680 21732 35736 21788
rect 35736 21732 35740 21788
rect 35676 21728 35740 21732
rect 35756 21788 35820 21792
rect 35756 21732 35760 21788
rect 35760 21732 35816 21788
rect 35816 21732 35820 21788
rect 35756 21728 35820 21732
rect 35836 21788 35900 21792
rect 35836 21732 35840 21788
rect 35840 21732 35896 21788
rect 35896 21732 35900 21788
rect 35836 21728 35900 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 4876 20700 4940 20704
rect 4876 20644 4880 20700
rect 4880 20644 4936 20700
rect 4936 20644 4940 20700
rect 4876 20640 4940 20644
rect 4956 20700 5020 20704
rect 4956 20644 4960 20700
rect 4960 20644 5016 20700
rect 5016 20644 5020 20700
rect 4956 20640 5020 20644
rect 5036 20700 5100 20704
rect 5036 20644 5040 20700
rect 5040 20644 5096 20700
rect 5096 20644 5100 20700
rect 5036 20640 5100 20644
rect 5116 20700 5180 20704
rect 5116 20644 5120 20700
rect 5120 20644 5176 20700
rect 5176 20644 5180 20700
rect 5116 20640 5180 20644
rect 35596 20700 35660 20704
rect 35596 20644 35600 20700
rect 35600 20644 35656 20700
rect 35656 20644 35660 20700
rect 35596 20640 35660 20644
rect 35676 20700 35740 20704
rect 35676 20644 35680 20700
rect 35680 20644 35736 20700
rect 35736 20644 35740 20700
rect 35676 20640 35740 20644
rect 35756 20700 35820 20704
rect 35756 20644 35760 20700
rect 35760 20644 35816 20700
rect 35816 20644 35820 20700
rect 35756 20640 35820 20644
rect 35836 20700 35900 20704
rect 35836 20644 35840 20700
rect 35840 20644 35896 20700
rect 35896 20644 35900 20700
rect 35836 20640 35900 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 4876 19612 4940 19616
rect 4876 19556 4880 19612
rect 4880 19556 4936 19612
rect 4936 19556 4940 19612
rect 4876 19552 4940 19556
rect 4956 19612 5020 19616
rect 4956 19556 4960 19612
rect 4960 19556 5016 19612
rect 5016 19556 5020 19612
rect 4956 19552 5020 19556
rect 5036 19612 5100 19616
rect 5036 19556 5040 19612
rect 5040 19556 5096 19612
rect 5096 19556 5100 19612
rect 5036 19552 5100 19556
rect 5116 19612 5180 19616
rect 5116 19556 5120 19612
rect 5120 19556 5176 19612
rect 5176 19556 5180 19612
rect 5116 19552 5180 19556
rect 35596 19612 35660 19616
rect 35596 19556 35600 19612
rect 35600 19556 35656 19612
rect 35656 19556 35660 19612
rect 35596 19552 35660 19556
rect 35676 19612 35740 19616
rect 35676 19556 35680 19612
rect 35680 19556 35736 19612
rect 35736 19556 35740 19612
rect 35676 19552 35740 19556
rect 35756 19612 35820 19616
rect 35756 19556 35760 19612
rect 35760 19556 35816 19612
rect 35816 19556 35820 19612
rect 35756 19552 35820 19556
rect 35836 19612 35900 19616
rect 35836 19556 35840 19612
rect 35840 19556 35896 19612
rect 35896 19556 35900 19612
rect 35836 19552 35900 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 4876 18524 4940 18528
rect 4876 18468 4880 18524
rect 4880 18468 4936 18524
rect 4936 18468 4940 18524
rect 4876 18464 4940 18468
rect 4956 18524 5020 18528
rect 4956 18468 4960 18524
rect 4960 18468 5016 18524
rect 5016 18468 5020 18524
rect 4956 18464 5020 18468
rect 5036 18524 5100 18528
rect 5036 18468 5040 18524
rect 5040 18468 5096 18524
rect 5096 18468 5100 18524
rect 5036 18464 5100 18468
rect 5116 18524 5180 18528
rect 5116 18468 5120 18524
rect 5120 18468 5176 18524
rect 5176 18468 5180 18524
rect 5116 18464 5180 18468
rect 35596 18524 35660 18528
rect 35596 18468 35600 18524
rect 35600 18468 35656 18524
rect 35656 18468 35660 18524
rect 35596 18464 35660 18468
rect 35676 18524 35740 18528
rect 35676 18468 35680 18524
rect 35680 18468 35736 18524
rect 35736 18468 35740 18524
rect 35676 18464 35740 18468
rect 35756 18524 35820 18528
rect 35756 18468 35760 18524
rect 35760 18468 35816 18524
rect 35816 18468 35820 18524
rect 35756 18464 35820 18468
rect 35836 18524 35900 18528
rect 35836 18468 35840 18524
rect 35840 18468 35896 18524
rect 35896 18468 35900 18524
rect 35836 18464 35900 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 4876 17436 4940 17440
rect 4876 17380 4880 17436
rect 4880 17380 4936 17436
rect 4936 17380 4940 17436
rect 4876 17376 4940 17380
rect 4956 17436 5020 17440
rect 4956 17380 4960 17436
rect 4960 17380 5016 17436
rect 5016 17380 5020 17436
rect 4956 17376 5020 17380
rect 5036 17436 5100 17440
rect 5036 17380 5040 17436
rect 5040 17380 5096 17436
rect 5096 17380 5100 17436
rect 5036 17376 5100 17380
rect 5116 17436 5180 17440
rect 5116 17380 5120 17436
rect 5120 17380 5176 17436
rect 5176 17380 5180 17436
rect 5116 17376 5180 17380
rect 35596 17436 35660 17440
rect 35596 17380 35600 17436
rect 35600 17380 35656 17436
rect 35656 17380 35660 17436
rect 35596 17376 35660 17380
rect 35676 17436 35740 17440
rect 35676 17380 35680 17436
rect 35680 17380 35736 17436
rect 35736 17380 35740 17436
rect 35676 17376 35740 17380
rect 35756 17436 35820 17440
rect 35756 17380 35760 17436
rect 35760 17380 35816 17436
rect 35816 17380 35820 17436
rect 35756 17376 35820 17380
rect 35836 17436 35900 17440
rect 35836 17380 35840 17436
rect 35840 17380 35896 17436
rect 35896 17380 35900 17436
rect 35836 17376 35900 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 4876 16348 4940 16352
rect 4876 16292 4880 16348
rect 4880 16292 4936 16348
rect 4936 16292 4940 16348
rect 4876 16288 4940 16292
rect 4956 16348 5020 16352
rect 4956 16292 4960 16348
rect 4960 16292 5016 16348
rect 5016 16292 5020 16348
rect 4956 16288 5020 16292
rect 5036 16348 5100 16352
rect 5036 16292 5040 16348
rect 5040 16292 5096 16348
rect 5096 16292 5100 16348
rect 5036 16288 5100 16292
rect 5116 16348 5180 16352
rect 5116 16292 5120 16348
rect 5120 16292 5176 16348
rect 5176 16292 5180 16348
rect 5116 16288 5180 16292
rect 35596 16348 35660 16352
rect 35596 16292 35600 16348
rect 35600 16292 35656 16348
rect 35656 16292 35660 16348
rect 35596 16288 35660 16292
rect 35676 16348 35740 16352
rect 35676 16292 35680 16348
rect 35680 16292 35736 16348
rect 35736 16292 35740 16348
rect 35676 16288 35740 16292
rect 35756 16348 35820 16352
rect 35756 16292 35760 16348
rect 35760 16292 35816 16348
rect 35816 16292 35820 16348
rect 35756 16288 35820 16292
rect 35836 16348 35900 16352
rect 35836 16292 35840 16348
rect 35840 16292 35896 16348
rect 35896 16292 35900 16348
rect 35836 16288 35900 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 4876 15260 4940 15264
rect 4876 15204 4880 15260
rect 4880 15204 4936 15260
rect 4936 15204 4940 15260
rect 4876 15200 4940 15204
rect 4956 15260 5020 15264
rect 4956 15204 4960 15260
rect 4960 15204 5016 15260
rect 5016 15204 5020 15260
rect 4956 15200 5020 15204
rect 5036 15260 5100 15264
rect 5036 15204 5040 15260
rect 5040 15204 5096 15260
rect 5096 15204 5100 15260
rect 5036 15200 5100 15204
rect 5116 15260 5180 15264
rect 5116 15204 5120 15260
rect 5120 15204 5176 15260
rect 5176 15204 5180 15260
rect 5116 15200 5180 15204
rect 35596 15260 35660 15264
rect 35596 15204 35600 15260
rect 35600 15204 35656 15260
rect 35656 15204 35660 15260
rect 35596 15200 35660 15204
rect 35676 15260 35740 15264
rect 35676 15204 35680 15260
rect 35680 15204 35736 15260
rect 35736 15204 35740 15260
rect 35676 15200 35740 15204
rect 35756 15260 35820 15264
rect 35756 15204 35760 15260
rect 35760 15204 35816 15260
rect 35816 15204 35820 15260
rect 35756 15200 35820 15204
rect 35836 15260 35900 15264
rect 35836 15204 35840 15260
rect 35840 15204 35896 15260
rect 35896 15204 35900 15260
rect 35836 15200 35900 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 4876 14172 4940 14176
rect 4876 14116 4880 14172
rect 4880 14116 4936 14172
rect 4936 14116 4940 14172
rect 4876 14112 4940 14116
rect 4956 14172 5020 14176
rect 4956 14116 4960 14172
rect 4960 14116 5016 14172
rect 5016 14116 5020 14172
rect 4956 14112 5020 14116
rect 5036 14172 5100 14176
rect 5036 14116 5040 14172
rect 5040 14116 5096 14172
rect 5096 14116 5100 14172
rect 5036 14112 5100 14116
rect 5116 14172 5180 14176
rect 5116 14116 5120 14172
rect 5120 14116 5176 14172
rect 5176 14116 5180 14172
rect 5116 14112 5180 14116
rect 35596 14172 35660 14176
rect 35596 14116 35600 14172
rect 35600 14116 35656 14172
rect 35656 14116 35660 14172
rect 35596 14112 35660 14116
rect 35676 14172 35740 14176
rect 35676 14116 35680 14172
rect 35680 14116 35736 14172
rect 35736 14116 35740 14172
rect 35676 14112 35740 14116
rect 35756 14172 35820 14176
rect 35756 14116 35760 14172
rect 35760 14116 35816 14172
rect 35816 14116 35820 14172
rect 35756 14112 35820 14116
rect 35836 14172 35900 14176
rect 35836 14116 35840 14172
rect 35840 14116 35896 14172
rect 35896 14116 35900 14172
rect 35836 14112 35900 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 4876 13084 4940 13088
rect 4876 13028 4880 13084
rect 4880 13028 4936 13084
rect 4936 13028 4940 13084
rect 4876 13024 4940 13028
rect 4956 13084 5020 13088
rect 4956 13028 4960 13084
rect 4960 13028 5016 13084
rect 5016 13028 5020 13084
rect 4956 13024 5020 13028
rect 5036 13084 5100 13088
rect 5036 13028 5040 13084
rect 5040 13028 5096 13084
rect 5096 13028 5100 13084
rect 5036 13024 5100 13028
rect 5116 13084 5180 13088
rect 5116 13028 5120 13084
rect 5120 13028 5176 13084
rect 5176 13028 5180 13084
rect 5116 13024 5180 13028
rect 35596 13084 35660 13088
rect 35596 13028 35600 13084
rect 35600 13028 35656 13084
rect 35656 13028 35660 13084
rect 35596 13024 35660 13028
rect 35676 13084 35740 13088
rect 35676 13028 35680 13084
rect 35680 13028 35736 13084
rect 35736 13028 35740 13084
rect 35676 13024 35740 13028
rect 35756 13084 35820 13088
rect 35756 13028 35760 13084
rect 35760 13028 35816 13084
rect 35816 13028 35820 13084
rect 35756 13024 35820 13028
rect 35836 13084 35900 13088
rect 35836 13028 35840 13084
rect 35840 13028 35896 13084
rect 35896 13028 35900 13084
rect 35836 13024 35900 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 4876 11996 4940 12000
rect 4876 11940 4880 11996
rect 4880 11940 4936 11996
rect 4936 11940 4940 11996
rect 4876 11936 4940 11940
rect 4956 11996 5020 12000
rect 4956 11940 4960 11996
rect 4960 11940 5016 11996
rect 5016 11940 5020 11996
rect 4956 11936 5020 11940
rect 5036 11996 5100 12000
rect 5036 11940 5040 11996
rect 5040 11940 5096 11996
rect 5096 11940 5100 11996
rect 5036 11936 5100 11940
rect 5116 11996 5180 12000
rect 5116 11940 5120 11996
rect 5120 11940 5176 11996
rect 5176 11940 5180 11996
rect 5116 11936 5180 11940
rect 35596 11996 35660 12000
rect 35596 11940 35600 11996
rect 35600 11940 35656 11996
rect 35656 11940 35660 11996
rect 35596 11936 35660 11940
rect 35676 11996 35740 12000
rect 35676 11940 35680 11996
rect 35680 11940 35736 11996
rect 35736 11940 35740 11996
rect 35676 11936 35740 11940
rect 35756 11996 35820 12000
rect 35756 11940 35760 11996
rect 35760 11940 35816 11996
rect 35816 11940 35820 11996
rect 35756 11936 35820 11940
rect 35836 11996 35900 12000
rect 35836 11940 35840 11996
rect 35840 11940 35896 11996
rect 35896 11940 35900 11996
rect 35836 11936 35900 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 4876 10908 4940 10912
rect 4876 10852 4880 10908
rect 4880 10852 4936 10908
rect 4936 10852 4940 10908
rect 4876 10848 4940 10852
rect 4956 10908 5020 10912
rect 4956 10852 4960 10908
rect 4960 10852 5016 10908
rect 5016 10852 5020 10908
rect 4956 10848 5020 10852
rect 5036 10908 5100 10912
rect 5036 10852 5040 10908
rect 5040 10852 5096 10908
rect 5096 10852 5100 10908
rect 5036 10848 5100 10852
rect 5116 10908 5180 10912
rect 5116 10852 5120 10908
rect 5120 10852 5176 10908
rect 5176 10852 5180 10908
rect 5116 10848 5180 10852
rect 35596 10908 35660 10912
rect 35596 10852 35600 10908
rect 35600 10852 35656 10908
rect 35656 10852 35660 10908
rect 35596 10848 35660 10852
rect 35676 10908 35740 10912
rect 35676 10852 35680 10908
rect 35680 10852 35736 10908
rect 35736 10852 35740 10908
rect 35676 10848 35740 10852
rect 35756 10908 35820 10912
rect 35756 10852 35760 10908
rect 35760 10852 35816 10908
rect 35816 10852 35820 10908
rect 35756 10848 35820 10852
rect 35836 10908 35900 10912
rect 35836 10852 35840 10908
rect 35840 10852 35896 10908
rect 35896 10852 35900 10908
rect 35836 10848 35900 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 4876 9820 4940 9824
rect 4876 9764 4880 9820
rect 4880 9764 4936 9820
rect 4936 9764 4940 9820
rect 4876 9760 4940 9764
rect 4956 9820 5020 9824
rect 4956 9764 4960 9820
rect 4960 9764 5016 9820
rect 5016 9764 5020 9820
rect 4956 9760 5020 9764
rect 5036 9820 5100 9824
rect 5036 9764 5040 9820
rect 5040 9764 5096 9820
rect 5096 9764 5100 9820
rect 5036 9760 5100 9764
rect 5116 9820 5180 9824
rect 5116 9764 5120 9820
rect 5120 9764 5176 9820
rect 5176 9764 5180 9820
rect 5116 9760 5180 9764
rect 35596 9820 35660 9824
rect 35596 9764 35600 9820
rect 35600 9764 35656 9820
rect 35656 9764 35660 9820
rect 35596 9760 35660 9764
rect 35676 9820 35740 9824
rect 35676 9764 35680 9820
rect 35680 9764 35736 9820
rect 35736 9764 35740 9820
rect 35676 9760 35740 9764
rect 35756 9820 35820 9824
rect 35756 9764 35760 9820
rect 35760 9764 35816 9820
rect 35816 9764 35820 9820
rect 35756 9760 35820 9764
rect 35836 9820 35900 9824
rect 35836 9764 35840 9820
rect 35840 9764 35896 9820
rect 35896 9764 35900 9820
rect 35836 9760 35900 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 4876 8732 4940 8736
rect 4876 8676 4880 8732
rect 4880 8676 4936 8732
rect 4936 8676 4940 8732
rect 4876 8672 4940 8676
rect 4956 8732 5020 8736
rect 4956 8676 4960 8732
rect 4960 8676 5016 8732
rect 5016 8676 5020 8732
rect 4956 8672 5020 8676
rect 5036 8732 5100 8736
rect 5036 8676 5040 8732
rect 5040 8676 5096 8732
rect 5096 8676 5100 8732
rect 5036 8672 5100 8676
rect 5116 8732 5180 8736
rect 5116 8676 5120 8732
rect 5120 8676 5176 8732
rect 5176 8676 5180 8732
rect 5116 8672 5180 8676
rect 35596 8732 35660 8736
rect 35596 8676 35600 8732
rect 35600 8676 35656 8732
rect 35656 8676 35660 8732
rect 35596 8672 35660 8676
rect 35676 8732 35740 8736
rect 35676 8676 35680 8732
rect 35680 8676 35736 8732
rect 35736 8676 35740 8732
rect 35676 8672 35740 8676
rect 35756 8732 35820 8736
rect 35756 8676 35760 8732
rect 35760 8676 35816 8732
rect 35816 8676 35820 8732
rect 35756 8672 35820 8676
rect 35836 8732 35900 8736
rect 35836 8676 35840 8732
rect 35840 8676 35896 8732
rect 35896 8676 35900 8732
rect 35836 8672 35900 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 35596 7644 35660 7648
rect 35596 7588 35600 7644
rect 35600 7588 35656 7644
rect 35656 7588 35660 7644
rect 35596 7584 35660 7588
rect 35676 7644 35740 7648
rect 35676 7588 35680 7644
rect 35680 7588 35736 7644
rect 35736 7588 35740 7644
rect 35676 7584 35740 7588
rect 35756 7644 35820 7648
rect 35756 7588 35760 7644
rect 35760 7588 35816 7644
rect 35816 7588 35820 7644
rect 35756 7584 35820 7588
rect 35836 7644 35900 7648
rect 35836 7588 35840 7644
rect 35840 7588 35896 7644
rect 35896 7588 35900 7644
rect 35836 7584 35900 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 35596 6556 35660 6560
rect 35596 6500 35600 6556
rect 35600 6500 35656 6556
rect 35656 6500 35660 6556
rect 35596 6496 35660 6500
rect 35676 6556 35740 6560
rect 35676 6500 35680 6556
rect 35680 6500 35736 6556
rect 35736 6500 35740 6556
rect 35676 6496 35740 6500
rect 35756 6556 35820 6560
rect 35756 6500 35760 6556
rect 35760 6500 35816 6556
rect 35816 6500 35820 6556
rect 35756 6496 35820 6500
rect 35836 6556 35900 6560
rect 35836 6500 35840 6556
rect 35840 6500 35896 6556
rect 35896 6500 35900 6556
rect 35836 6496 35900 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 35596 5468 35660 5472
rect 35596 5412 35600 5468
rect 35600 5412 35656 5468
rect 35656 5412 35660 5468
rect 35596 5408 35660 5412
rect 35676 5468 35740 5472
rect 35676 5412 35680 5468
rect 35680 5412 35736 5468
rect 35736 5412 35740 5468
rect 35676 5408 35740 5412
rect 35756 5468 35820 5472
rect 35756 5412 35760 5468
rect 35760 5412 35816 5468
rect 35816 5412 35820 5468
rect 35756 5408 35820 5412
rect 35836 5468 35900 5472
rect 35836 5412 35840 5468
rect 35840 5412 35896 5468
rect 35896 5412 35900 5468
rect 35836 5408 35900 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 35596 4380 35660 4384
rect 35596 4324 35600 4380
rect 35600 4324 35656 4380
rect 35656 4324 35660 4380
rect 35596 4320 35660 4324
rect 35676 4380 35740 4384
rect 35676 4324 35680 4380
rect 35680 4324 35736 4380
rect 35736 4324 35740 4380
rect 35676 4320 35740 4324
rect 35756 4380 35820 4384
rect 35756 4324 35760 4380
rect 35760 4324 35816 4380
rect 35816 4324 35820 4380
rect 35756 4320 35820 4324
rect 35836 4380 35900 4384
rect 35836 4324 35840 4380
rect 35840 4324 35896 4380
rect 35896 4324 35900 4380
rect 35836 4320 35900 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 35596 3292 35660 3296
rect 35596 3236 35600 3292
rect 35600 3236 35656 3292
rect 35656 3236 35660 3292
rect 35596 3232 35660 3236
rect 35676 3292 35740 3296
rect 35676 3236 35680 3292
rect 35680 3236 35736 3292
rect 35736 3236 35740 3292
rect 35676 3232 35740 3236
rect 35756 3292 35820 3296
rect 35756 3236 35760 3292
rect 35760 3236 35816 3292
rect 35816 3236 35820 3292
rect 35756 3232 35820 3236
rect 35836 3292 35900 3296
rect 35836 3236 35840 3292
rect 35840 3236 35896 3292
rect 35896 3236 35900 3292
rect 35836 3232 35900 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
rect 35596 2204 35660 2208
rect 35596 2148 35600 2204
rect 35600 2148 35656 2204
rect 35656 2148 35660 2204
rect 35596 2144 35660 2148
rect 35676 2204 35740 2208
rect 35676 2148 35680 2204
rect 35680 2148 35736 2204
rect 35736 2148 35740 2204
rect 35676 2144 35740 2148
rect 35756 2204 35820 2208
rect 35756 2148 35760 2204
rect 35760 2148 35816 2204
rect 35816 2148 35820 2204
rect 35756 2144 35820 2148
rect 35836 2204 35900 2208
rect 35836 2148 35840 2204
rect 35840 2148 35896 2204
rect 35896 2148 35900 2204
rect 35836 2144 35900 2148
<< metal4 >>
rect 4208 38656 4528 38672
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 36260 4528 36416
rect 4208 36024 4250 36260
rect 4486 36024 4528 36260
rect 4208 35392 4528 36024
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5624 4528 5952
rect 4208 5388 4250 5624
rect 4486 5388 4528 5624
rect 4208 4928 4528 5388
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 38112 5188 38672
rect 4868 38048 4876 38112
rect 4940 38048 4956 38112
rect 5020 38048 5036 38112
rect 5100 38048 5116 38112
rect 5180 38048 5188 38112
rect 4868 37024 5188 38048
rect 4868 36960 4876 37024
rect 4940 36960 4956 37024
rect 5020 36960 5036 37024
rect 5100 36960 5116 37024
rect 5180 36960 5188 37024
rect 4868 36920 5188 36960
rect 4868 36684 4910 36920
rect 5146 36684 5188 36920
rect 4868 35936 5188 36684
rect 4868 35872 4876 35936
rect 4940 35872 4956 35936
rect 5020 35872 5036 35936
rect 5100 35872 5116 35936
rect 5180 35872 5188 35936
rect 4868 34848 5188 35872
rect 4868 34784 4876 34848
rect 4940 34784 4956 34848
rect 5020 34784 5036 34848
rect 5100 34784 5116 34848
rect 5180 34784 5188 34848
rect 4868 33760 5188 34784
rect 4868 33696 4876 33760
rect 4940 33696 4956 33760
rect 5020 33696 5036 33760
rect 5100 33696 5116 33760
rect 5180 33696 5188 33760
rect 4868 32672 5188 33696
rect 4868 32608 4876 32672
rect 4940 32608 4956 32672
rect 5020 32608 5036 32672
rect 5100 32608 5116 32672
rect 5180 32608 5188 32672
rect 4868 31584 5188 32608
rect 4868 31520 4876 31584
rect 4940 31520 4956 31584
rect 5020 31520 5036 31584
rect 5100 31520 5116 31584
rect 5180 31520 5188 31584
rect 4868 30496 5188 31520
rect 4868 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5188 30496
rect 4868 29408 5188 30432
rect 4868 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5188 29408
rect 4868 28320 5188 29344
rect 4868 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5188 28320
rect 4868 27232 5188 28256
rect 4868 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5188 27232
rect 4868 26144 5188 27168
rect 4868 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5188 26144
rect 4868 25056 5188 26080
rect 4868 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5188 25056
rect 4868 23968 5188 24992
rect 4868 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5188 23968
rect 4868 22880 5188 23904
rect 4868 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5188 22880
rect 4868 21792 5188 22816
rect 4868 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5188 21792
rect 4868 20704 5188 21728
rect 4868 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5188 20704
rect 4868 19616 5188 20640
rect 4868 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5188 19616
rect 4868 18528 5188 19552
rect 4868 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5188 18528
rect 4868 17440 5188 18464
rect 4868 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5188 17440
rect 4868 16352 5188 17376
rect 4868 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5188 16352
rect 4868 15264 5188 16288
rect 4868 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5188 15264
rect 4868 14176 5188 15200
rect 4868 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5188 14176
rect 4868 13088 5188 14112
rect 4868 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5188 13088
rect 4868 12000 5188 13024
rect 4868 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5188 12000
rect 4868 10912 5188 11936
rect 4868 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5188 10912
rect 4868 9824 5188 10848
rect 4868 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5188 9824
rect 4868 8736 5188 9760
rect 4868 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5188 8736
rect 4868 7648 5188 8672
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 6284 5188 6496
rect 4868 6048 4910 6284
rect 5146 6048 5188 6284
rect 4868 5472 5188 6048
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
rect 34928 38656 35248 38672
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 36260 35248 36416
rect 34928 36024 34970 36260
rect 35206 36024 35248 36260
rect 34928 35392 35248 36024
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 5624 35248 5952
rect 34928 5388 34970 5624
rect 35206 5388 35248 5624
rect 34928 4928 35248 5388
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
rect 35588 38112 35908 38672
rect 35588 38048 35596 38112
rect 35660 38048 35676 38112
rect 35740 38048 35756 38112
rect 35820 38048 35836 38112
rect 35900 38048 35908 38112
rect 35588 37024 35908 38048
rect 35588 36960 35596 37024
rect 35660 36960 35676 37024
rect 35740 36960 35756 37024
rect 35820 36960 35836 37024
rect 35900 36960 35908 37024
rect 35588 36920 35908 36960
rect 35588 36684 35630 36920
rect 35866 36684 35908 36920
rect 35588 35936 35908 36684
rect 35588 35872 35596 35936
rect 35660 35872 35676 35936
rect 35740 35872 35756 35936
rect 35820 35872 35836 35936
rect 35900 35872 35908 35936
rect 35588 34848 35908 35872
rect 35588 34784 35596 34848
rect 35660 34784 35676 34848
rect 35740 34784 35756 34848
rect 35820 34784 35836 34848
rect 35900 34784 35908 34848
rect 35588 33760 35908 34784
rect 35588 33696 35596 33760
rect 35660 33696 35676 33760
rect 35740 33696 35756 33760
rect 35820 33696 35836 33760
rect 35900 33696 35908 33760
rect 35588 32672 35908 33696
rect 35588 32608 35596 32672
rect 35660 32608 35676 32672
rect 35740 32608 35756 32672
rect 35820 32608 35836 32672
rect 35900 32608 35908 32672
rect 35588 31584 35908 32608
rect 35588 31520 35596 31584
rect 35660 31520 35676 31584
rect 35740 31520 35756 31584
rect 35820 31520 35836 31584
rect 35900 31520 35908 31584
rect 35588 30496 35908 31520
rect 35588 30432 35596 30496
rect 35660 30432 35676 30496
rect 35740 30432 35756 30496
rect 35820 30432 35836 30496
rect 35900 30432 35908 30496
rect 35588 29408 35908 30432
rect 35588 29344 35596 29408
rect 35660 29344 35676 29408
rect 35740 29344 35756 29408
rect 35820 29344 35836 29408
rect 35900 29344 35908 29408
rect 35588 28320 35908 29344
rect 35588 28256 35596 28320
rect 35660 28256 35676 28320
rect 35740 28256 35756 28320
rect 35820 28256 35836 28320
rect 35900 28256 35908 28320
rect 35588 27232 35908 28256
rect 35588 27168 35596 27232
rect 35660 27168 35676 27232
rect 35740 27168 35756 27232
rect 35820 27168 35836 27232
rect 35900 27168 35908 27232
rect 35588 26144 35908 27168
rect 35588 26080 35596 26144
rect 35660 26080 35676 26144
rect 35740 26080 35756 26144
rect 35820 26080 35836 26144
rect 35900 26080 35908 26144
rect 35588 25056 35908 26080
rect 35588 24992 35596 25056
rect 35660 24992 35676 25056
rect 35740 24992 35756 25056
rect 35820 24992 35836 25056
rect 35900 24992 35908 25056
rect 35588 23968 35908 24992
rect 35588 23904 35596 23968
rect 35660 23904 35676 23968
rect 35740 23904 35756 23968
rect 35820 23904 35836 23968
rect 35900 23904 35908 23968
rect 35588 22880 35908 23904
rect 35588 22816 35596 22880
rect 35660 22816 35676 22880
rect 35740 22816 35756 22880
rect 35820 22816 35836 22880
rect 35900 22816 35908 22880
rect 35588 21792 35908 22816
rect 35588 21728 35596 21792
rect 35660 21728 35676 21792
rect 35740 21728 35756 21792
rect 35820 21728 35836 21792
rect 35900 21728 35908 21792
rect 35588 20704 35908 21728
rect 35588 20640 35596 20704
rect 35660 20640 35676 20704
rect 35740 20640 35756 20704
rect 35820 20640 35836 20704
rect 35900 20640 35908 20704
rect 35588 19616 35908 20640
rect 35588 19552 35596 19616
rect 35660 19552 35676 19616
rect 35740 19552 35756 19616
rect 35820 19552 35836 19616
rect 35900 19552 35908 19616
rect 35588 18528 35908 19552
rect 35588 18464 35596 18528
rect 35660 18464 35676 18528
rect 35740 18464 35756 18528
rect 35820 18464 35836 18528
rect 35900 18464 35908 18528
rect 35588 17440 35908 18464
rect 35588 17376 35596 17440
rect 35660 17376 35676 17440
rect 35740 17376 35756 17440
rect 35820 17376 35836 17440
rect 35900 17376 35908 17440
rect 35588 16352 35908 17376
rect 35588 16288 35596 16352
rect 35660 16288 35676 16352
rect 35740 16288 35756 16352
rect 35820 16288 35836 16352
rect 35900 16288 35908 16352
rect 35588 15264 35908 16288
rect 35588 15200 35596 15264
rect 35660 15200 35676 15264
rect 35740 15200 35756 15264
rect 35820 15200 35836 15264
rect 35900 15200 35908 15264
rect 35588 14176 35908 15200
rect 35588 14112 35596 14176
rect 35660 14112 35676 14176
rect 35740 14112 35756 14176
rect 35820 14112 35836 14176
rect 35900 14112 35908 14176
rect 35588 13088 35908 14112
rect 35588 13024 35596 13088
rect 35660 13024 35676 13088
rect 35740 13024 35756 13088
rect 35820 13024 35836 13088
rect 35900 13024 35908 13088
rect 35588 12000 35908 13024
rect 35588 11936 35596 12000
rect 35660 11936 35676 12000
rect 35740 11936 35756 12000
rect 35820 11936 35836 12000
rect 35900 11936 35908 12000
rect 35588 10912 35908 11936
rect 35588 10848 35596 10912
rect 35660 10848 35676 10912
rect 35740 10848 35756 10912
rect 35820 10848 35836 10912
rect 35900 10848 35908 10912
rect 35588 9824 35908 10848
rect 35588 9760 35596 9824
rect 35660 9760 35676 9824
rect 35740 9760 35756 9824
rect 35820 9760 35836 9824
rect 35900 9760 35908 9824
rect 35588 8736 35908 9760
rect 35588 8672 35596 8736
rect 35660 8672 35676 8736
rect 35740 8672 35756 8736
rect 35820 8672 35836 8736
rect 35900 8672 35908 8736
rect 35588 7648 35908 8672
rect 35588 7584 35596 7648
rect 35660 7584 35676 7648
rect 35740 7584 35756 7648
rect 35820 7584 35836 7648
rect 35900 7584 35908 7648
rect 35588 6560 35908 7584
rect 35588 6496 35596 6560
rect 35660 6496 35676 6560
rect 35740 6496 35756 6560
rect 35820 6496 35836 6560
rect 35900 6496 35908 6560
rect 35588 6284 35908 6496
rect 35588 6048 35630 6284
rect 35866 6048 35908 6284
rect 35588 5472 35908 6048
rect 35588 5408 35596 5472
rect 35660 5408 35676 5472
rect 35740 5408 35756 5472
rect 35820 5408 35836 5472
rect 35900 5408 35908 5472
rect 35588 4384 35908 5408
rect 35588 4320 35596 4384
rect 35660 4320 35676 4384
rect 35740 4320 35756 4384
rect 35820 4320 35836 4384
rect 35900 4320 35908 4384
rect 35588 3296 35908 4320
rect 35588 3232 35596 3296
rect 35660 3232 35676 3296
rect 35740 3232 35756 3296
rect 35820 3232 35836 3296
rect 35900 3232 35908 3296
rect 35588 2208 35908 3232
rect 35588 2144 35596 2208
rect 35660 2144 35676 2208
rect 35740 2144 35756 2208
rect 35820 2144 35836 2208
rect 35900 2144 35908 2208
rect 35588 2128 35908 2144
<< via4 >>
rect 4250 36024 4486 36260
rect 4250 5388 4486 5624
rect 4910 36684 5146 36920
rect 4910 6048 5146 6284
rect 34970 36024 35206 36260
rect 34970 5388 35206 5624
rect 35630 36684 35866 36920
rect 35630 6048 35866 6284
<< metal5 >>
rect 1056 36920 37676 36962
rect 1056 36684 4910 36920
rect 5146 36684 35630 36920
rect 35866 36684 37676 36920
rect 1056 36642 37676 36684
rect 1056 36260 37676 36302
rect 1056 36024 4250 36260
rect 4486 36024 34970 36260
rect 35206 36024 37676 36260
rect 1056 35982 37676 36024
rect 1056 6284 37676 6326
rect 1056 6048 4910 6284
rect 5146 6048 35630 6284
rect 35866 6048 37676 6284
rect 1056 6006 37676 6048
rect 1056 5624 37676 5666
rect 1056 5388 4250 5624
rect 4486 5388 34970 5624
rect 35206 5388 37676 5624
rect 1056 5346 37676 5388
use sky130_fd_sc_hd__fill_2  FILLER_0_3 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1668240031
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1668240031
transform 1 0 1840 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1668240031
transform 1 0 2944 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1668240031
transform 1 0 3772 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1668240031
transform 1 0 4140 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37
timestamp 1668240031
transform 1 0 4508 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1668240031
transform 1 0 5612 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55
timestamp 1668240031
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57
timestamp 1668240031
transform 1 0 6348 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63
timestamp 1668240031
transform 1 0 6900 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67
timestamp 1668240031
transform 1 0 7268 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_79
timestamp 1668240031
transform 1 0 8372 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83
timestamp 1668240031
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_85
timestamp 1668240031
transform 1 0 8924 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_96
timestamp 1668240031
transform 1 0 9936 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_103
timestamp 1668240031
transform 1 0 10580 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1668240031
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 1668240031
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_135
timestamp 1668240031
transform 1 0 13524 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_139
timestamp 1668240031
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_141
timestamp 1668240031
transform 1 0 14076 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_152
timestamp 1668240031
transform 1 0 15088 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_159
timestamp 1668240031
transform 1 0 15732 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1668240031
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_169
timestamp 1668240031
transform 1 0 16652 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_186
timestamp 1668240031
transform 1 0 18216 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1668240031
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1668240031
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_202
timestamp 1668240031
transform 1 0 19688 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_215
timestamp 1668240031
transform 1 0 20884 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1668240031
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1668240031
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_230
timestamp 1668240031
transform 1 0 22264 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_245
timestamp 1668240031
transform 1 0 23644 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_251
timestamp 1668240031
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1668240031
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_258
timestamp 1668240031
transform 1 0 24840 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_265
timestamp 1668240031
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 1668240031
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_281
timestamp 1668240031
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_293
timestamp 1668240031
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp 1668240031
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 1668240031
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_317
timestamp 1668240031
transform 1 0 30268 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_329
timestamp 1668240031
transform 1 0 31372 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_335
timestamp 1668240031
transform 1 0 31924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 1668240031
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_349
timestamp 1668240031
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp 1668240031
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_365
timestamp 1668240031
transform 1 0 34684 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_370
timestamp 1668240031
transform 1 0 35144 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_382
timestamp 1668240031
transform 1 0 36248 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_386
timestamp 1668240031
transform 1 0 36616 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_390
timestamp 1668240031
transform 1 0 36984 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_393
timestamp 1668240031
transform 1 0 37260 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1668240031
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_8
timestamp 1668240031
transform 1 0 1840 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_20
timestamp 1668240031
transform 1 0 2944 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_32
timestamp 1668240031
transform 1 0 4048 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_44
timestamp 1668240031
transform 1 0 5152 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1668240031
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1668240031
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1668240031
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1668240031
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_105
timestamp 1668240031
transform 1 0 10764 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1668240031
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_113
timestamp 1668240031
transform 1 0 11500 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_118
timestamp 1668240031
transform 1 0 11960 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_142
timestamp 1668240031
transform 1 0 14168 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_166
timestamp 1668240031
transform 1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_169
timestamp 1668240031
transform 1 0 16652 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_173
timestamp 1668240031
transform 1 0 17020 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_194
timestamp 1668240031
transform 1 0 18952 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_205
timestamp 1668240031
transform 1 0 19964 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_218
timestamp 1668240031
transform 1 0 21160 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_1_225
timestamp 1668240031
transform 1 0 21804 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_237
timestamp 1668240031
transform 1 0 22908 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1668240031
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1668240031
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1668240031
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1668240031
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1668240031
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_305
timestamp 1668240031
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_317
timestamp 1668240031
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1668240031
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1668240031
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1668240031
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1668240031
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_361
timestamp 1668240031
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_373
timestamp 1668240031
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_385
timestamp 1668240031
transform 1 0 36524 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_390
timestamp 1668240031
transform 1 0 36984 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_393
timestamp 1668240031
transform 1 0 37260 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1668240031
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1668240031
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1668240031
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1668240031
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1668240031
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1668240031
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1668240031
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1668240031
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1668240031
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_85
timestamp 1668240031
transform 1 0 8924 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_93
timestamp 1668240031
transform 1 0 9660 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_98
timestamp 1668240031
transform 1 0 10120 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_122
timestamp 1668240031
transform 1 0 12328 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_135
timestamp 1668240031
transform 1 0 13524 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1668240031
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_141
timestamp 1668240031
transform 1 0 14076 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_147
timestamp 1668240031
transform 1 0 14628 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_157
timestamp 1668240031
transform 1 0 15548 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_174
timestamp 1668240031
transform 1 0 17112 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_181
timestamp 1668240031
transform 1 0 17756 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_194
timestamp 1668240031
transform 1 0 18952 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_197
timestamp 1668240031
transform 1 0 19228 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_205
timestamp 1668240031
transform 1 0 19964 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_228
timestamp 1668240031
transform 1 0 22080 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_241
timestamp 1668240031
transform 1 0 23276 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_248
timestamp 1668240031
transform 1 0 23920 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_253
timestamp 1668240031
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_258
timestamp 1668240031
transform 1 0 24840 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_270
timestamp 1668240031
transform 1 0 25944 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_282
timestamp 1668240031
transform 1 0 27048 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_290
timestamp 1668240031
transform 1 0 27784 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_295
timestamp 1668240031
transform 1 0 28244 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_305
timestamp 1668240031
transform 1 0 29164 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1668240031
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1668240031
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1668240031
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1668240031
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1668240031
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1668240031
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1668240031
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1668240031
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_389
timestamp 1668240031
transform 1 0 36892 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_393
timestamp 1668240031
transform 1 0 37260 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1668240031
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1668240031
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1668240031
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1668240031
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1668240031
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1668240031
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1668240031
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1668240031
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1668240031
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_93
timestamp 1668240031
transform 1 0 9660 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_110
timestamp 1668240031
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_113
timestamp 1668240031
transform 1 0 11500 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_119
timestamp 1668240031
transform 1 0 12052 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_129
timestamp 1668240031
transform 1 0 12972 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_142
timestamp 1668240031
transform 1 0 14168 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_166
timestamp 1668240031
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_169
timestamp 1668240031
transform 1 0 16652 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_173
timestamp 1668240031
transform 1 0 17020 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_194
timestamp 1668240031
transform 1 0 18952 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_218
timestamp 1668240031
transform 1 0 21160 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_225
timestamp 1668240031
transform 1 0 21804 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_247
timestamp 1668240031
transform 1 0 23828 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_260
timestamp 1668240031
transform 1 0 25024 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_272
timestamp 1668240031
transform 1 0 26128 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_281
timestamp 1668240031
transform 1 0 26956 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_304
timestamp 1668240031
transform 1 0 29072 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_317
timestamp 1668240031
transform 1 0 30268 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_324
timestamp 1668240031
transform 1 0 30912 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1668240031
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1668240031
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1668240031
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1668240031
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1668240031
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1668240031
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_393
timestamp 1668240031
transform 1 0 37260 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1668240031
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1668240031
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1668240031
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1668240031
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1668240031
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1668240031
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1668240031
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1668240031
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1668240031
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1668240031
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_97
timestamp 1668240031
transform 1 0 10028 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_103
timestamp 1668240031
transform 1 0 10580 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_116
timestamp 1668240031
transform 1 0 11776 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_129
timestamp 1668240031
transform 1 0 12972 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_138
timestamp 1668240031
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_141
timestamp 1668240031
transform 1 0 14076 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_152
timestamp 1668240031
transform 1 0 15088 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_160
timestamp 1668240031
transform 1 0 15824 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_170
timestamp 1668240031
transform 1 0 16744 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_180
timestamp 1668240031
transform 1 0 17664 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_193
timestamp 1668240031
transform 1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_197
timestamp 1668240031
transform 1 0 19228 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_206
timestamp 1668240031
transform 1 0 20056 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_213
timestamp 1668240031
transform 1 0 20700 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_228
timestamp 1668240031
transform 1 0 22080 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_241
timestamp 1668240031
transform 1 0 23276 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_249
timestamp 1668240031
transform 1 0 24012 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1668240031
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1668240031
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_277
timestamp 1668240031
transform 1 0 26588 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_285
timestamp 1668240031
transform 1 0 27324 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_290
timestamp 1668240031
transform 1 0 27784 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_303
timestamp 1668240031
transform 1 0 28980 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1668240031
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_309
timestamp 1668240031
transform 1 0 29532 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_331
timestamp 1668240031
transform 1 0 31556 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_338
timestamp 1668240031
transform 1 0 32200 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1668240031
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1668240031
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1668240031
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1668240031
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1668240031
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_389
timestamp 1668240031
transform 1 0 36892 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_393
timestamp 1668240031
transform 1 0 37260 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1668240031
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1668240031
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1668240031
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1668240031
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1668240031
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1668240031
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1668240031
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1668240031
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1668240031
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_93
timestamp 1668240031
transform 1 0 9660 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_99
timestamp 1668240031
transform 1 0 10212 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_103
timestamp 1668240031
transform 1 0 10580 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_110
timestamp 1668240031
transform 1 0 11224 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_113
timestamp 1668240031
transform 1 0 11500 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_117
timestamp 1668240031
transform 1 0 11868 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_121
timestamp 1668240031
transform 1 0 12236 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_134
timestamp 1668240031
transform 1 0 13432 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_158
timestamp 1668240031
transform 1 0 15640 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_5_165
timestamp 1668240031
transform 1 0 16284 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_169
timestamp 1668240031
transform 1 0 16652 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_174
timestamp 1668240031
transform 1 0 17112 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_189
timestamp 1668240031
transform 1 0 18492 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_201
timestamp 1668240031
transform 1 0 19596 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_213
timestamp 1668240031
transform 1 0 20700 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_221
timestamp 1668240031
transform 1 0 21436 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1668240031
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1668240031
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1668240031
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1668240031
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1668240031
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1668240031
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_281
timestamp 1668240031
transform 1 0 26956 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_293
timestamp 1668240031
transform 1 0 28060 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_297
timestamp 1668240031
transform 1 0 28428 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_301
timestamp 1668240031
transform 1 0 28796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_314
timestamp 1668240031
transform 1 0 29992 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_327
timestamp 1668240031
transform 1 0 31188 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_334
timestamp 1668240031
transform 1 0 31832 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_337
timestamp 1668240031
transform 1 0 32108 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_348
timestamp 1668240031
transform 1 0 33120 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_357
timestamp 1668240031
transform 1 0 33948 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_369
timestamp 1668240031
transform 1 0 35052 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_381
timestamp 1668240031
transform 1 0 36156 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_389
timestamp 1668240031
transform 1 0 36892 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_393
timestamp 1668240031
transform 1 0 37260 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1668240031
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_8
timestamp 1668240031
transform 1 0 1840 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_20
timestamp 1668240031
transform 1 0 2944 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1668240031
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1668240031
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1668240031
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1668240031
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1668240031
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1668240031
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1668240031
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1668240031
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_109
timestamp 1668240031
transform 1 0 11132 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_131
timestamp 1668240031
transform 1 0 13156 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_138
timestamp 1668240031
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_141
timestamp 1668240031
transform 1 0 14076 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_152
timestamp 1668240031
transform 1 0 15088 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_6_180
timestamp 1668240031
transform 1 0 17664 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_192
timestamp 1668240031
transform 1 0 18768 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1668240031
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1668240031
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1668240031
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1668240031
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1668240031
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1668240031
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1668240031
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_265
timestamp 1668240031
transform 1 0 25484 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_6_291
timestamp 1668240031
transform 1 0 27876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_306
timestamp 1668240031
transform 1 0 29256 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_309
timestamp 1668240031
transform 1 0 29532 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_313
timestamp 1668240031
transform 1 0 29900 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_317
timestamp 1668240031
transform 1 0 30268 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_323
timestamp 1668240031
transform 1 0 30820 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_344
timestamp 1668240031
transform 1 0 32752 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1668240031
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1668240031
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1668240031
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1668240031
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_392
timestamp 1668240031
transform 1 0 37168 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1668240031
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1668240031
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1668240031
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1668240031
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1668240031
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1668240031
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1668240031
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1668240031
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1668240031
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1668240031
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1668240031
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1668240031
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_113
timestamp 1668240031
transform 1 0 11500 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_7_119
timestamp 1668240031
transform 1 0 12052 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_7_134
timestamp 1668240031
transform 1 0 13432 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_142
timestamp 1668240031
transform 1 0 14168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_152
timestamp 1668240031
transform 1 0 15088 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_7_165
timestamp 1668240031
transform 1 0 16284 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_169
timestamp 1668240031
transform 1 0 16652 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_174
timestamp 1668240031
transform 1 0 17112 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_186
timestamp 1668240031
transform 1 0 18216 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_198
timestamp 1668240031
transform 1 0 19320 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_210
timestamp 1668240031
transform 1 0 20424 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_222
timestamp 1668240031
transform 1 0 21528 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1668240031
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1668240031
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1668240031
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1668240031
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_273
timestamp 1668240031
transform 1 0 26220 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_278
timestamp 1668240031
transform 1 0 26680 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_281
timestamp 1668240031
transform 1 0 26956 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_292
timestamp 1668240031
transform 1 0 27968 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_299
timestamp 1668240031
transform 1 0 28612 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_323
timestamp 1668240031
transform 1 0 30820 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_330
timestamp 1668240031
transform 1 0 31464 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_7_337
timestamp 1668240031
transform 1 0 32108 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_363
timestamp 1668240031
transform 1 0 34500 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_370
timestamp 1668240031
transform 1 0 35144 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_382
timestamp 1668240031
transform 1 0 36248 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_390
timestamp 1668240031
transform 1 0 36984 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_393
timestamp 1668240031
transform 1 0 37260 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1668240031
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1668240031
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1668240031
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1668240031
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1668240031
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1668240031
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1668240031
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1668240031
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1668240031
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1668240031
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1668240031
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_109
timestamp 1668240031
transform 1 0 11132 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_115
timestamp 1668240031
transform 1 0 11684 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_136
timestamp 1668240031
transform 1 0 13616 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1668240031
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_153
timestamp 1668240031
transform 1 0 15180 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_165
timestamp 1668240031
transform 1 0 16284 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_172
timestamp 1668240031
transform 1 0 16928 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_184
timestamp 1668240031
transform 1 0 18032 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1668240031
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1668240031
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1668240031
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1668240031
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1668240031
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1668240031
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1668240031
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_265
timestamp 1668240031
transform 1 0 25484 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_293
timestamp 1668240031
transform 1 0 28060 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_306
timestamp 1668240031
transform 1 0 29256 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_309
timestamp 1668240031
transform 1 0 29532 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_320
timestamp 1668240031
transform 1 0 30544 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_333
timestamp 1668240031
transform 1 0 31740 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_346
timestamp 1668240031
transform 1 0 32936 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_353
timestamp 1668240031
transform 1 0 33580 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_360
timestamp 1668240031
transform 1 0 34224 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1668240031
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1668240031
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_389
timestamp 1668240031
transform 1 0 36892 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_393
timestamp 1668240031
transform 1 0 37260 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1668240031
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1668240031
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1668240031
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1668240031
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1668240031
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1668240031
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1668240031
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_89
timestamp 1668240031
transform 1 0 9292 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_101
timestamp 1668240031
transform 1 0 10396 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_109
timestamp 1668240031
transform 1 0 11132 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_113
timestamp 1668240031
transform 1 0 11500 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_119
timestamp 1668240031
transform 1 0 12052 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_123
timestamp 1668240031
transform 1 0 12420 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_130
timestamp 1668240031
transform 1 0 13064 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_134
timestamp 1668240031
transform 1 0 13432 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_155
timestamp 1668240031
transform 1 0 15364 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_162
timestamp 1668240031
transform 1 0 16008 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1668240031
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1668240031
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1668240031
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1668240031
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1668240031
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1668240031
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1668240031
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1668240031
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_249
timestamp 1668240031
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_261
timestamp 1668240031
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1668240031
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1668240031
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_281
timestamp 1668240031
transform 1 0 26956 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_286
timestamp 1668240031
transform 1 0 27416 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_293
timestamp 1668240031
transform 1 0 28060 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_301
timestamp 1668240031
transform 1 0 28796 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_323
timestamp 1668240031
transform 1 0 30820 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_330
timestamp 1668240031
transform 1 0 31464 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_9_337
timestamp 1668240031
transform 1 0 32108 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_343
timestamp 1668240031
transform 1 0 32660 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_364
timestamp 1668240031
transform 1 0 34592 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_376
timestamp 1668240031
transform 1 0 35696 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_388
timestamp 1668240031
transform 1 0 36800 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_393
timestamp 1668240031
transform 1 0 37260 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1668240031
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1668240031
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1668240031
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1668240031
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1668240031
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_53
timestamp 1668240031
transform 1 0 5980 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_70
timestamp 1668240031
transform 1 0 7544 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1668240031
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1668240031
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_85
timestamp 1668240031
transform 1 0 8924 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_90
timestamp 1668240031
transform 1 0 9384 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_102
timestamp 1668240031
transform 1 0 10488 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_106
timestamp 1668240031
transform 1 0 10856 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_118
timestamp 1668240031
transform 1 0 11960 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_126
timestamp 1668240031
transform 1 0 12696 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_138
timestamp 1668240031
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_141
timestamp 1668240031
transform 1 0 14076 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_146
timestamp 1668240031
transform 1 0 14536 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_161
timestamp 1668240031
transform 1 0 15916 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_168
timestamp 1668240031
transform 1 0 16560 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_174
timestamp 1668240031
transform 1 0 17112 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_178
timestamp 1668240031
transform 1 0 17480 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_190
timestamp 1668240031
transform 1 0 18584 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1668240031
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1668240031
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1668240031
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1668240031
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1668240031
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1668240031
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_253
timestamp 1668240031
transform 1 0 24380 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_261
timestamp 1668240031
transform 1 0 25116 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_266
timestamp 1668240031
transform 1 0 25576 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_278
timestamp 1668240031
transform 1 0 26680 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_282
timestamp 1668240031
transform 1 0 27048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_286
timestamp 1668240031
transform 1 0 27416 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_294
timestamp 1668240031
transform 1 0 28152 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_305
timestamp 1668240031
transform 1 0 29164 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_309
timestamp 1668240031
transform 1 0 29532 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_320
timestamp 1668240031
transform 1 0 30544 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_324
timestamp 1668240031
transform 1 0 30912 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_345
timestamp 1668240031
transform 1 0 32844 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_358
timestamp 1668240031
transform 1 0 34040 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_365
timestamp 1668240031
transform 1 0 34684 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_370
timestamp 1668240031
transform 1 0 35144 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_382
timestamp 1668240031
transform 1 0 36248 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1668240031
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1668240031
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1668240031
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1668240031
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp 1668240031
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_57
timestamp 1668240031
transform 1 0 6348 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_79
timestamp 1668240031
transform 1 0 8372 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_87
timestamp 1668240031
transform 1 0 9108 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp 1668240031
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_113
timestamp 1668240031
transform 1 0 11500 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_117
timestamp 1668240031
transform 1 0 11868 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_121
timestamp 1668240031
transform 1 0 12236 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_133
timestamp 1668240031
transform 1 0 13340 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_137
timestamp 1668240031
transform 1 0 13708 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_150
timestamp 1668240031
transform 1 0 14904 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_11_165
timestamp 1668240031
transform 1 0 16284 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_169
timestamp 1668240031
transform 1 0 16652 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_191
timestamp 1668240031
transform 1 0 18676 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_203
timestamp 1668240031
transform 1 0 19780 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_215
timestamp 1668240031
transform 1 0 20884 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1668240031
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1668240031
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1668240031
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_249
timestamp 1668240031
transform 1 0 24012 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_257
timestamp 1668240031
transform 1 0 24748 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_271
timestamp 1668240031
transform 1 0 26036 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_278
timestamp 1668240031
transform 1 0 26680 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_281
timestamp 1668240031
transform 1 0 26956 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_296
timestamp 1668240031
transform 1 0 28336 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_320
timestamp 1668240031
transform 1 0 30544 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_327
timestamp 1668240031
transform 1 0 31188 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_334
timestamp 1668240031
transform 1 0 31832 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_337
timestamp 1668240031
transform 1 0 32108 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_348
timestamp 1668240031
transform 1 0 33120 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_361
timestamp 1668240031
transform 1 0 34316 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_368
timestamp 1668240031
transform 1 0 34960 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_380
timestamp 1668240031
transform 1 0 36064 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_393
timestamp 1668240031
transform 1 0 37260 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1668240031
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1668240031
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1668240031
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1668240031
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1668240031
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_56
timestamp 1668240031
transform 1 0 6256 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_69
timestamp 1668240031
transform 1 0 7452 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_82
timestamp 1668240031
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_85
timestamp 1668240031
transform 1 0 8924 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_100
timestamp 1668240031
transform 1 0 10304 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_107
timestamp 1668240031
transform 1 0 10948 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_114
timestamp 1668240031
transform 1 0 11592 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_118
timestamp 1668240031
transform 1 0 11960 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_128
timestamp 1668240031
transform 1 0 12880 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_134
timestamp 1668240031
transform 1 0 13432 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_138
timestamp 1668240031
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_141
timestamp 1668240031
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_163
timestamp 1668240031
transform 1 0 16100 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_175
timestamp 1668240031
transform 1 0 17204 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_187
timestamp 1668240031
transform 1 0 18308 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1668240031
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1668240031
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1668240031
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1668240031
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_233
timestamp 1668240031
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1668240031
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1668240031
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_253
timestamp 1668240031
transform 1 0 24380 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_276
timestamp 1668240031
transform 1 0 26496 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_300
timestamp 1668240031
transform 1 0 28704 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_309
timestamp 1668240031
transform 1 0 29532 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_322
timestamp 1668240031
transform 1 0 30728 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_328
timestamp 1668240031
transform 1 0 31280 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_338
timestamp 1668240031
transform 1 0 32200 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_351
timestamp 1668240031
transform 1 0 33396 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_355
timestamp 1668240031
transform 1 0 33764 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_359
timestamp 1668240031
transform 1 0 34132 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1668240031
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1668240031
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1668240031
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_389
timestamp 1668240031
transform 1 0 36892 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_393
timestamp 1668240031
transform 1 0 37260 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 1668240031
transform 1 0 1380 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_8
timestamp 1668240031
transform 1 0 1840 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_20
timestamp 1668240031
transform 1 0 2944 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_32
timestamp 1668240031
transform 1 0 4048 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_44
timestamp 1668240031
transform 1 0 5152 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_57
timestamp 1668240031
transform 1 0 6348 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_63
timestamp 1668240031
transform 1 0 6900 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_73
timestamp 1668240031
transform 1 0 7820 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_79
timestamp 1668240031
transform 1 0 8372 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_89
timestamp 1668240031
transform 1 0 9292 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_102
timestamp 1668240031
transform 1 0 10488 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_106
timestamp 1668240031
transform 1 0 10856 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_110
timestamp 1668240031
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_113
timestamp 1668240031
transform 1 0 11500 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_135
timestamp 1668240031
transform 1 0 13524 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_148
timestamp 1668240031
transform 1 0 14720 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_160
timestamp 1668240031
transform 1 0 15824 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1668240031
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1668240031
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1668240031
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_205
timestamp 1668240031
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1668240031
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1668240031
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_225
timestamp 1668240031
transform 1 0 21804 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_233
timestamp 1668240031
transform 1 0 22540 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_240
timestamp 1668240031
transform 1 0 23184 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_244
timestamp 1668240031
transform 1 0 23552 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_248
timestamp 1668240031
transform 1 0 23920 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_256
timestamp 1668240031
transform 1 0 24656 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_260
timestamp 1668240031
transform 1 0 25024 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_267
timestamp 1668240031
transform 1 0 25668 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_274
timestamp 1668240031
transform 1 0 26312 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_281
timestamp 1668240031
transform 1 0 26956 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_292
timestamp 1668240031
transform 1 0 27968 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_305
timestamp 1668240031
transform 1 0 29164 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_313
timestamp 1668240031
transform 1 0 29900 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_334
timestamp 1668240031
transform 1 0 31832 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_337
timestamp 1668240031
transform 1 0 32108 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_13_365
timestamp 1668240031
transform 1 0 34684 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_377
timestamp 1668240031
transform 1 0 35788 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_385
timestamp 1668240031
transform 1 0 36524 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_390
timestamp 1668240031
transform 1 0 36984 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_393
timestamp 1668240031
transform 1 0 37260 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1668240031
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1668240031
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1668240031
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1668240031
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1668240031
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_53
timestamp 1668240031
transform 1 0 5980 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_74
timestamp 1668240031
transform 1 0 7912 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_78
timestamp 1668240031
transform 1 0 8280 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1668240031
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_85
timestamp 1668240031
transform 1 0 8924 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_107
timestamp 1668240031
transform 1 0 10948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_113
timestamp 1668240031
transform 1 0 11500 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_117
timestamp 1668240031
transform 1 0 11868 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_130
timestamp 1668240031
transform 1 0 13064 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_138
timestamp 1668240031
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1668240031
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1668240031
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1668240031
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1668240031
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1668240031
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1668240031
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1668240031
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1668240031
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_221
timestamp 1668240031
transform 1 0 21436 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_229
timestamp 1668240031
transform 1 0 22172 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_250
timestamp 1668240031
transform 1 0 24104 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_253
timestamp 1668240031
transform 1 0 24380 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_275
timestamp 1668240031
transform 1 0 26404 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_298
timestamp 1668240031
transform 1 0 28520 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_305
timestamp 1668240031
transform 1 0 29164 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_309
timestamp 1668240031
transform 1 0 29532 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_320
timestamp 1668240031
transform 1 0 30544 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_330
timestamp 1668240031
transform 1 0 31464 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_336
timestamp 1668240031
transform 1 0 32016 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_346
timestamp 1668240031
transform 1 0 32936 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_353
timestamp 1668240031
transform 1 0 33580 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_360
timestamp 1668240031
transform 1 0 34224 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1668240031
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1668240031
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_389
timestamp 1668240031
transform 1 0 36892 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_393
timestamp 1668240031
transform 1 0 37260 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1668240031
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1668240031
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1668240031
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1668240031
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1668240031
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1668240031
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_57
timestamp 1668240031
transform 1 0 6348 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_68
timestamp 1668240031
transform 1 0 7360 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_75
timestamp 1668240031
transform 1 0 8004 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_79
timestamp 1668240031
transform 1 0 8372 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_100
timestamp 1668240031
transform 1 0 10304 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_107
timestamp 1668240031
transform 1 0 10948 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1668240031
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_113
timestamp 1668240031
transform 1 0 11500 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_119
timestamp 1668240031
transform 1 0 12052 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_141
timestamp 1668240031
transform 1 0 14076 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_153
timestamp 1668240031
transform 1 0 15180 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_165
timestamp 1668240031
transform 1 0 16284 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_169
timestamp 1668240031
transform 1 0 16652 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_15_183
timestamp 1668240031
transform 1 0 17940 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_195
timestamp 1668240031
transform 1 0 19044 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_207
timestamp 1668240031
transform 1 0 20148 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_219
timestamp 1668240031
transform 1 0 21252 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1668240031
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_225
timestamp 1668240031
transform 1 0 21804 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_236
timestamp 1668240031
transform 1 0 22816 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_246
timestamp 1668240031
transform 1 0 23736 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_254
timestamp 1668240031
transform 1 0 24472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_261
timestamp 1668240031
transform 1 0 25116 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_274
timestamp 1668240031
transform 1 0 26312 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_15_281
timestamp 1668240031
transform 1 0 26956 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_289
timestamp 1668240031
transform 1 0 27692 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_313
timestamp 1668240031
transform 1 0 29900 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_326
timestamp 1668240031
transform 1 0 31096 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_333
timestamp 1668240031
transform 1 0 31740 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_337
timestamp 1668240031
transform 1 0 32108 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_342
timestamp 1668240031
transform 1 0 32568 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_355
timestamp 1668240031
transform 1 0 33764 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_362
timestamp 1668240031
transform 1 0 34408 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_374
timestamp 1668240031
transform 1 0 35512 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_386
timestamp 1668240031
transform 1 0 36616 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_393
timestamp 1668240031
transform 1 0 37260 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1668240031
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1668240031
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1668240031
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1668240031
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1668240031
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_53
timestamp 1668240031
transform 1 0 5980 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_60
timestamp 1668240031
transform 1 0 6624 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_68
timestamp 1668240031
transform 1 0 7360 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_74
timestamp 1668240031
transform 1 0 7912 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1668240031
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_85
timestamp 1668240031
transform 1 0 8924 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_94
timestamp 1668240031
transform 1 0 9752 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_118
timestamp 1668240031
transform 1 0 11960 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_131
timestamp 1668240031
transform 1 0 13156 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1668240031
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1668240031
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1668240031
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1668240031
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_177
timestamp 1668240031
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1668240031
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1668240031
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1668240031
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_209
timestamp 1668240031
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_221
timestamp 1668240031
transform 1 0 21436 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_229
timestamp 1668240031
transform 1 0 22172 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_233
timestamp 1668240031
transform 1 0 22540 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_240
timestamp 1668240031
transform 1 0 23184 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_246
timestamp 1668240031
transform 1 0 23736 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_250
timestamp 1668240031
transform 1 0 24104 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_253
timestamp 1668240031
transform 1 0 24380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_264
timestamp 1668240031
transform 1 0 25392 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_272
timestamp 1668240031
transform 1 0 26128 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_282
timestamp 1668240031
transform 1 0 27048 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_295
timestamp 1668240031
transform 1 0 28244 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_305
timestamp 1668240031
transform 1 0 29164 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_309
timestamp 1668240031
transform 1 0 29532 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_332
timestamp 1668240031
transform 1 0 31648 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_356
timestamp 1668240031
transform 1 0 33856 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_365
timestamp 1668240031
transform 1 0 34684 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_370
timestamp 1668240031
transform 1 0 35144 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_382
timestamp 1668240031
transform 1 0 36248 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1668240031
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1668240031
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1668240031
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1668240031
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1668240031
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1668240031
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_57
timestamp 1668240031
transform 1 0 6348 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_68
timestamp 1668240031
transform 1 0 7360 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_75
timestamp 1668240031
transform 1 0 8004 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_82
timestamp 1668240031
transform 1 0 8648 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_95
timestamp 1668240031
transform 1 0 9844 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp 1668240031
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_113
timestamp 1668240031
transform 1 0 11500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_126
timestamp 1668240031
transform 1 0 12696 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_17_140
timestamp 1668240031
transform 1 0 13984 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_152
timestamp 1668240031
transform 1 0 15088 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_164
timestamp 1668240031
transform 1 0 16192 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1668240031
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 1668240031
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_193
timestamp 1668240031
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_205
timestamp 1668240031
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1668240031
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1668240031
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_225
timestamp 1668240031
transform 1 0 21804 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_247
timestamp 1668240031
transform 1 0 23828 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_260
timestamp 1668240031
transform 1 0 25024 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1668240031
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1668240031
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_281
timestamp 1668240031
transform 1 0 26956 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_292
timestamp 1668240031
transform 1 0 27968 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_299
timestamp 1668240031
transform 1 0 28612 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_306
timestamp 1668240031
transform 1 0 29256 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_310
timestamp 1668240031
transform 1 0 29624 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_320
timestamp 1668240031
transform 1 0 30544 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_324
timestamp 1668240031
transform 1 0 30912 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_334
timestamp 1668240031
transform 1 0 31832 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_337
timestamp 1668240031
transform 1 0 32108 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_342
timestamp 1668240031
transform 1 0 32568 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_346
timestamp 1668240031
transform 1 0 32936 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_367
timestamp 1668240031
transform 1 0 34868 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_379
timestamp 1668240031
transform 1 0 35972 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1668240031
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_393
timestamp 1668240031
transform 1 0 37260 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1668240031
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1668240031
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1668240031
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1668240031
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1668240031
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_53
timestamp 1668240031
transform 1 0 5980 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_58
timestamp 1668240031
transform 1 0 6440 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1668240031
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_85
timestamp 1668240031
transform 1 0 8924 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_96
timestamp 1668240031
transform 1 0 9936 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_105
timestamp 1668240031
transform 1 0 10764 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_112
timestamp 1668240031
transform 1 0 11408 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_136
timestamp 1668240031
transform 1 0 13616 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_141
timestamp 1668240031
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_146
timestamp 1668240031
transform 1 0 14536 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_158
timestamp 1668240031
transform 1 0 15640 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_170
timestamp 1668240031
transform 1 0 16744 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_182
timestamp 1668240031
transform 1 0 17848 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1668240031
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_197
timestamp 1668240031
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_209
timestamp 1668240031
transform 1 0 20332 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_237
timestamp 1668240031
transform 1 0 22908 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_250
timestamp 1668240031
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_253
timestamp 1668240031
transform 1 0 24380 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_279
timestamp 1668240031
transform 1 0 26772 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_303
timestamp 1668240031
transform 1 0 28980 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1668240031
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_309
timestamp 1668240031
transform 1 0 29532 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_314
timestamp 1668240031
transform 1 0 29992 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_321
timestamp 1668240031
transform 1 0 30636 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_329
timestamp 1668240031
transform 1 0 31372 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_340
timestamp 1668240031
transform 1 0 32384 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_353
timestamp 1668240031
transform 1 0 33580 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_360
timestamp 1668240031
transform 1 0 34224 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_365
timestamp 1668240031
transform 1 0 34684 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_370
timestamp 1668240031
transform 1 0 35144 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_382
timestamp 1668240031
transform 1 0 36248 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1668240031
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1668240031
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1668240031
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1668240031
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1668240031
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1668240031
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_57
timestamp 1668240031
transform 1 0 6348 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_79
timestamp 1668240031
transform 1 0 8372 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_96
timestamp 1668240031
transform 1 0 9936 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_100
timestamp 1668240031
transform 1 0 10304 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_110
timestamp 1668240031
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_113
timestamp 1668240031
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_124
timestamp 1668240031
transform 1 0 12512 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_138
timestamp 1668240031
transform 1 0 13800 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_145
timestamp 1668240031
transform 1 0 14444 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_157
timestamp 1668240031
transform 1 0 15548 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_165
timestamp 1668240031
transform 1 0 16284 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_19_169
timestamp 1668240031
transform 1 0 16652 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_175
timestamp 1668240031
transform 1 0 17204 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_182
timestamp 1668240031
transform 1 0 17848 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_194
timestamp 1668240031
transform 1 0 18952 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_206
timestamp 1668240031
transform 1 0 20056 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_218
timestamp 1668240031
transform 1 0 21160 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_19_225
timestamp 1668240031
transform 1 0 21804 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_231
timestamp 1668240031
transform 1 0 22356 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_239
timestamp 1668240031
transform 1 0 23092 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_249
timestamp 1668240031
transform 1 0 24012 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_262
timestamp 1668240031
transform 1 0 25208 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_272
timestamp 1668240031
transform 1 0 26128 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_281
timestamp 1668240031
transform 1 0 26956 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_286
timestamp 1668240031
transform 1 0 27416 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_297
timestamp 1668240031
transform 1 0 28428 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_304
timestamp 1668240031
transform 1 0 29072 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_321
timestamp 1668240031
transform 1 0 30636 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_334
timestamp 1668240031
transform 1 0 31832 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_337
timestamp 1668240031
transform 1 0 32108 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_343
timestamp 1668240031
transform 1 0 32660 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_364
timestamp 1668240031
transform 1 0 34592 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_376
timestamp 1668240031
transform 1 0 35696 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_388
timestamp 1668240031
transform 1 0 36800 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_393
timestamp 1668240031
transform 1 0 37260 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1668240031
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_8
timestamp 1668240031
transform 1 0 1840 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_20
timestamp 1668240031
transform 1 0 2944 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1668240031
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1668240031
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_53
timestamp 1668240031
transform 1 0 5980 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_62
timestamp 1668240031
transform 1 0 6808 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_69
timestamp 1668240031
transform 1 0 7452 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_77
timestamp 1668240031
transform 1 0 8188 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_82
timestamp 1668240031
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_85
timestamp 1668240031
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_96
timestamp 1668240031
transform 1 0 9936 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_120
timestamp 1668240031
transform 1 0 12144 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_20_137
timestamp 1668240031
transform 1 0 13708 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_141
timestamp 1668240031
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_149
timestamp 1668240031
transform 1 0 14812 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_161
timestamp 1668240031
transform 1 0 15916 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_173
timestamp 1668240031
transform 1 0 17020 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_185
timestamp 1668240031
transform 1 0 18124 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_193
timestamp 1668240031
transform 1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1668240031
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_209
timestamp 1668240031
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_221
timestamp 1668240031
transform 1 0 21436 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_227
timestamp 1668240031
transform 1 0 21988 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_231
timestamp 1668240031
transform 1 0 22356 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_241
timestamp 1668240031
transform 1 0 23276 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_250
timestamp 1668240031
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_253
timestamp 1668240031
transform 1 0 24380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_264
timestamp 1668240031
transform 1 0 25392 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_274
timestamp 1668240031
transform 1 0 26312 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_20_302
timestamp 1668240031
transform 1 0 28888 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_309
timestamp 1668240031
transform 1 0 29532 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_331
timestamp 1668240031
transform 1 0 31556 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_355
timestamp 1668240031
transform 1 0 33764 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_362
timestamp 1668240031
transform 1 0 34408 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1668240031
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_377
timestamp 1668240031
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_392
timestamp 1668240031
transform 1 0 37168 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1668240031
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1668240031
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1668240031
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1668240031
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1668240031
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1668240031
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_57
timestamp 1668240031
transform 1 0 6348 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_63
timestamp 1668240031
transform 1 0 6900 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_73
timestamp 1668240031
transform 1 0 7820 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_77
timestamp 1668240031
transform 1 0 8188 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_98
timestamp 1668240031
transform 1 0 10120 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1668240031
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1668240031
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_113
timestamp 1668240031
transform 1 0 11500 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_139
timestamp 1668240031
transform 1 0 13892 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_146
timestamp 1668240031
transform 1 0 14536 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_158
timestamp 1668240031
transform 1 0 15640 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1668240031
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1668240031
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_181
timestamp 1668240031
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_193
timestamp 1668240031
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_205
timestamp 1668240031
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_217
timestamp 1668240031
transform 1 0 21068 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_222
timestamp 1668240031
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_225
timestamp 1668240031
transform 1 0 21804 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_237
timestamp 1668240031
transform 1 0 22908 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_250
timestamp 1668240031
transform 1 0 24104 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_278
timestamp 1668240031
transform 1 0 26680 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_281
timestamp 1668240031
transform 1 0 26956 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_290
timestamp 1668240031
transform 1 0 27784 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_305
timestamp 1668240031
transform 1 0 29164 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_312
timestamp 1668240031
transform 1 0 29808 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_319
timestamp 1668240031
transform 1 0 30452 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_326
timestamp 1668240031
transform 1 0 31096 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_21_333
timestamp 1668240031
transform 1 0 31740 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_337
timestamp 1668240031
transform 1 0 32108 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_350
timestamp 1668240031
transform 1 0 33304 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_354
timestamp 1668240031
transform 1 0 33672 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_358
timestamp 1668240031
transform 1 0 34040 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_370
timestamp 1668240031
transform 1 0 35144 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_382
timestamp 1668240031
transform 1 0 36248 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_390
timestamp 1668240031
transform 1 0 36984 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_393
timestamp 1668240031
transform 1 0 37260 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1668240031
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1668240031
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1668240031
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1668240031
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_41
timestamp 1668240031
transform 1 0 4876 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_50
timestamp 1668240031
transform 1 0 5704 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_74
timestamp 1668240031
transform 1 0 7912 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_78
timestamp 1668240031
transform 1 0 8280 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1668240031
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_85
timestamp 1668240031
transform 1 0 8924 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_98
timestamp 1668240031
transform 1 0 10120 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_111
timestamp 1668240031
transform 1 0 11316 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_124
timestamp 1668240031
transform 1 0 12512 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_136
timestamp 1668240031
transform 1 0 13616 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1668240031
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1668240031
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 1668240031
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_177
timestamp 1668240031
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1668240031
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1668240031
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1668240031
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_209
timestamp 1668240031
transform 1 0 20332 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_217
timestamp 1668240031
transform 1 0 21068 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_238
timestamp 1668240031
transform 1 0 23000 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1668240031
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1668240031
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_253
timestamp 1668240031
transform 1 0 24380 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_279
timestamp 1668240031
transform 1 0 26772 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_290
timestamp 1668240031
transform 1 0 27784 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1668240031
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1668240031
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_309
timestamp 1668240031
transform 1 0 29532 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_319
timestamp 1668240031
transform 1 0 30452 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_326
timestamp 1668240031
transform 1 0 31096 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_333
timestamp 1668240031
transform 1 0 31740 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_337
timestamp 1668240031
transform 1 0 32108 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_341
timestamp 1668240031
transform 1 0 32476 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_348
timestamp 1668240031
transform 1 0 33120 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_356
timestamp 1668240031
transform 1 0 33856 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_361
timestamp 1668240031
transform 1 0 34316 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_365
timestamp 1668240031
transform 1 0 34684 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_376
timestamp 1668240031
transform 1 0 35696 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_388
timestamp 1668240031
transform 1 0 36800 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1668240031
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1668240031
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1668240031
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1668240031
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_54
timestamp 1668240031
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_57
timestamp 1668240031
transform 1 0 6348 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_69
timestamp 1668240031
transform 1 0 7452 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_77
timestamp 1668240031
transform 1 0 8188 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_81
timestamp 1668240031
transform 1 0 8556 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1668240031
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1668240031
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_113
timestamp 1668240031
transform 1 0 11500 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_118
timestamp 1668240031
transform 1 0 11960 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_128
timestamp 1668240031
transform 1 0 12880 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_132
timestamp 1668240031
transform 1 0 13248 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_139
timestamp 1668240031
transform 1 0 13892 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_149
timestamp 1668240031
transform 1 0 14812 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_156
timestamp 1668240031
transform 1 0 15456 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1668240031
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_181
timestamp 1668240031
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_193
timestamp 1668240031
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_205
timestamp 1668240031
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1668240031
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1668240031
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_225
timestamp 1668240031
transform 1 0 21804 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_236
timestamp 1668240031
transform 1 0 22816 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_251
timestamp 1668240031
transform 1 0 24196 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_258
timestamp 1668240031
transform 1 0 24840 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_266
timestamp 1668240031
transform 1 0 25576 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_278
timestamp 1668240031
transform 1 0 26680 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_281
timestamp 1668240031
transform 1 0 26956 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_292
timestamp 1668240031
transform 1 0 27968 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_299
timestamp 1668240031
transform 1 0 28612 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_23_313
timestamp 1668240031
transform 1 0 29900 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_321
timestamp 1668240031
transform 1 0 30636 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_327
timestamp 1668240031
transform 1 0 31188 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_334
timestamp 1668240031
transform 1 0 31832 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_337
timestamp 1668240031
transform 1 0 32108 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_344
timestamp 1668240031
transform 1 0 32752 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_351
timestamp 1668240031
transform 1 0 33396 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_355
timestamp 1668240031
transform 1 0 33764 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_376
timestamp 1668240031
transform 1 0 35696 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_383
timestamp 1668240031
transform 1 0 36340 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1668240031
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_393
timestamp 1668240031
transform 1 0 37260 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1668240031
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1668240031
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1668240031
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1668240031
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_41
timestamp 1668240031
transform 1 0 4876 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_52
timestamp 1668240031
transform 1 0 5888 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_76
timestamp 1668240031
transform 1 0 8096 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_85
timestamp 1668240031
transform 1 0 8924 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_96
timestamp 1668240031
transform 1 0 9936 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_103
timestamp 1668240031
transform 1 0 10580 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_109
timestamp 1668240031
transform 1 0 11132 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_130
timestamp 1668240031
transform 1 0 13064 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1668240031
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_141
timestamp 1668240031
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_149
timestamp 1668240031
transform 1 0 14812 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_156
timestamp 1668240031
transform 1 0 15456 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_166
timestamp 1668240031
transform 1 0 16376 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_178
timestamp 1668240031
transform 1 0 17480 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_190
timestamp 1668240031
transform 1 0 18584 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1668240031
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_209
timestamp 1668240031
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_221
timestamp 1668240031
transform 1 0 21436 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_243
timestamp 1668240031
transform 1 0 23460 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1668240031
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_253
timestamp 1668240031
transform 1 0 24380 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_262
timestamp 1668240031
transform 1 0 25208 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_286
timestamp 1668240031
transform 1 0 27416 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_293
timestamp 1668240031
transform 1 0 28060 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_306
timestamp 1668240031
transform 1 0 29256 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_309
timestamp 1668240031
transform 1 0 29532 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_314
timestamp 1668240031
transform 1 0 29992 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_338
timestamp 1668240031
transform 1 0 32200 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_362
timestamp 1668240031
transform 1 0 34408 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_365
timestamp 1668240031
transform 1 0 34684 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_371
timestamp 1668240031
transform 1 0 35236 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_392
timestamp 1668240031
transform 1 0 37168 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1668240031
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1668240031
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1668240031
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1668240031
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1668240031
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1668240031
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_57
timestamp 1668240031
transform 1 0 6348 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_68
timestamp 1668240031
transform 1 0 7360 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_77
timestamp 1668240031
transform 1 0 8188 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_90
timestamp 1668240031
transform 1 0 9384 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_25_101
timestamp 1668240031
transform 1 0 10396 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_110
timestamp 1668240031
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_113
timestamp 1668240031
transform 1 0 11500 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_124
timestamp 1668240031
transform 1 0 12512 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_152
timestamp 1668240031
transform 1 0 15088 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_156
timestamp 1668240031
transform 1 0 15456 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_160
timestamp 1668240031
transform 1 0 15824 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_169
timestamp 1668240031
transform 1 0 16652 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_175
timestamp 1668240031
transform 1 0 17204 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_25_186
timestamp 1668240031
transform 1 0 18216 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_192
timestamp 1668240031
transform 1 0 18768 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_196
timestamp 1668240031
transform 1 0 19136 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_200
timestamp 1668240031
transform 1 0 19504 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_204
timestamp 1668240031
transform 1 0 19872 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_211
timestamp 1668240031
transform 1 0 20516 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1668240031
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_225
timestamp 1668240031
transform 1 0 21804 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_232
timestamp 1668240031
transform 1 0 22448 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_247
timestamp 1668240031
transform 1 0 23828 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_260
timestamp 1668240031
transform 1 0 25024 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1668240031
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1668240031
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_281
timestamp 1668240031
transform 1 0 26956 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_286
timestamp 1668240031
transform 1 0 27416 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_294
timestamp 1668240031
transform 1 0 28152 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_304
timestamp 1668240031
transform 1 0 29072 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_315
timestamp 1668240031
transform 1 0 30084 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_324
timestamp 1668240031
transform 1 0 30912 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_331
timestamp 1668240031
transform 1 0 31556 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1668240031
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_337
timestamp 1668240031
transform 1 0 32108 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_344
timestamp 1668240031
transform 1 0 32752 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_359
timestamp 1668240031
transform 1 0 34132 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_368
timestamp 1668240031
transform 1 0 34960 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_375
timestamp 1668240031
transform 1 0 35604 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_382
timestamp 1668240031
transform 1 0 36248 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_25_389
timestamp 1668240031
transform 1 0 36892 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_393
timestamp 1668240031
transform 1 0 37260 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1668240031
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1668240031
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1668240031
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1668240031
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1668240031
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_53
timestamp 1668240031
transform 1 0 5980 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_66
timestamp 1668240031
transform 1 0 7176 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_79
timestamp 1668240031
transform 1 0 8372 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1668240031
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_85
timestamp 1668240031
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_107
timestamp 1668240031
transform 1 0 10948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_113
timestamp 1668240031
transform 1 0 11500 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_117
timestamp 1668240031
transform 1 0 11868 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_130
timestamp 1668240031
transform 1 0 13064 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_137
timestamp 1668240031
transform 1 0 13708 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_141
timestamp 1668240031
transform 1 0 14076 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_149
timestamp 1668240031
transform 1 0 14812 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_155
timestamp 1668240031
transform 1 0 15364 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_159
timestamp 1668240031
transform 1 0 15732 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_166
timestamp 1668240031
transform 1 0 16376 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_170
timestamp 1668240031
transform 1 0 16744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_191
timestamp 1668240031
transform 1 0 18676 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1668240031
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_197
timestamp 1668240031
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_219
timestamp 1668240031
transform 1 0 21252 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_227
timestamp 1668240031
transform 1 0 21988 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_231
timestamp 1668240031
transform 1 0 22356 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_237
timestamp 1668240031
transform 1 0 22908 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_247
timestamp 1668240031
transform 1 0 23828 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1668240031
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_253
timestamp 1668240031
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_261
timestamp 1668240031
transform 1 0 25116 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_285
timestamp 1668240031
transform 1 0 27324 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_292
timestamp 1668240031
transform 1 0 27968 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_296
timestamp 1668240031
transform 1 0 28336 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_300
timestamp 1668240031
transform 1 0 28704 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_309
timestamp 1668240031
transform 1 0 29532 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_318
timestamp 1668240031
transform 1 0 30360 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_327
timestamp 1668240031
transform 1 0 31188 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_334
timestamp 1668240031
transform 1 0 31832 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_340
timestamp 1668240031
transform 1 0 32384 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_344
timestamp 1668240031
transform 1 0 32752 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_351
timestamp 1668240031
transform 1 0 33396 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_358
timestamp 1668240031
transform 1 0 34040 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_365
timestamp 1668240031
transform 1 0 34684 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_372
timestamp 1668240031
transform 1 0 35328 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_26_381
timestamp 1668240031
transform 1 0 36156 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_392
timestamp 1668240031
transform 1 0 37168 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1668240031
transform 1 0 1380 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_8
timestamp 1668240031
transform 1 0 1840 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_20
timestamp 1668240031
transform 1 0 2944 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_32
timestamp 1668240031
transform 1 0 4048 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_44
timestamp 1668240031
transform 1 0 5152 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_50
timestamp 1668240031
transform 1 0 5704 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp 1668240031
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_57
timestamp 1668240031
transform 1 0 6348 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_79
timestamp 1668240031
transform 1 0 8372 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_92
timestamp 1668240031
transform 1 0 9568 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1668240031
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1668240031
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_113
timestamp 1668240031
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_124
timestamp 1668240031
transform 1 0 12512 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_137
timestamp 1668240031
transform 1 0 13708 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_145
timestamp 1668240031
transform 1 0 14444 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1668240031
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1668240031
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_180
timestamp 1668240031
transform 1 0 17664 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_188
timestamp 1668240031
transform 1 0 18400 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_198
timestamp 1668240031
transform 1 0 19320 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_222
timestamp 1668240031
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_225
timestamp 1668240031
transform 1 0 21804 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_247
timestamp 1668240031
transform 1 0 23828 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_260
timestamp 1668240031
transform 1 0 25024 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 1668240031
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1668240031
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_281
timestamp 1668240031
transform 1 0 26956 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_286
timestamp 1668240031
transform 1 0 27416 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_294
timestamp 1668240031
transform 1 0 28152 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_303
timestamp 1668240031
transform 1 0 28980 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_310
timestamp 1668240031
transform 1 0 29624 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_334
timestamp 1668240031
transform 1 0 31832 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_337
timestamp 1668240031
transform 1 0 32108 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_359
timestamp 1668240031
transform 1 0 34132 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_387
timestamp 1668240031
transform 1 0 36708 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1668240031
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_393
timestamp 1668240031
transform 1 0 37260 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1668240031
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1668240031
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1668240031
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1668240031
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_41
timestamp 1668240031
transform 1 0 4876 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_49
timestamp 1668240031
transform 1 0 5612 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_54
timestamp 1668240031
transform 1 0 6072 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_67
timestamp 1668240031
transform 1 0 7268 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_28_78
timestamp 1668240031
transform 1 0 8280 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_28_85
timestamp 1668240031
transform 1 0 8924 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_94
timestamp 1668240031
transform 1 0 9752 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_107
timestamp 1668240031
transform 1 0 10948 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_131
timestamp 1668240031
transform 1 0 13156 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1668240031
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_141
timestamp 1668240031
transform 1 0 14076 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_147
timestamp 1668240031
transform 1 0 14628 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_157
timestamp 1668240031
transform 1 0 15548 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_167
timestamp 1668240031
transform 1 0 16468 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_180
timestamp 1668240031
transform 1 0 17664 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_184
timestamp 1668240031
transform 1 0 18032 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp 1668240031
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_197
timestamp 1668240031
transform 1 0 19228 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_214
timestamp 1668240031
transform 1 0 20792 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_221
timestamp 1668240031
transform 1 0 21436 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_225
timestamp 1668240031
transform 1 0 21804 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_229
timestamp 1668240031
transform 1 0 22172 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_236
timestamp 1668240031
transform 1 0 22816 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_28_249
timestamp 1668240031
transform 1 0 24012 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_253
timestamp 1668240031
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_258
timestamp 1668240031
transform 1 0 24840 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_271
timestamp 1668240031
transform 1 0 26036 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_295
timestamp 1668240031
transform 1 0 28244 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_304
timestamp 1668240031
transform 1 0 29072 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_309
timestamp 1668240031
transform 1 0 29532 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_318
timestamp 1668240031
transform 1 0 30360 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_326
timestamp 1668240031
transform 1 0 31096 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_347
timestamp 1668240031
transform 1 0 33028 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_358
timestamp 1668240031
transform 1 0 34040 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_28_365
timestamp 1668240031
transform 1 0 34684 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_371
timestamp 1668240031
transform 1 0 35236 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_378
timestamp 1668240031
transform 1 0 35880 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_390
timestamp 1668240031
transform 1 0 36984 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1668240031
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1668240031
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1668240031
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1668240031
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_54
timestamp 1668240031
transform 1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_57
timestamp 1668240031
transform 1 0 6348 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_29_68
timestamp 1668240031
transform 1 0 7360 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_79
timestamp 1668240031
transform 1 0 8372 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_86
timestamp 1668240031
transform 1 0 9016 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_110
timestamp 1668240031
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_113
timestamp 1668240031
transform 1 0 11500 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_117
timestamp 1668240031
transform 1 0 11868 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_121
timestamp 1668240031
transform 1 0 12236 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_145
timestamp 1668240031
transform 1 0 14444 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_158
timestamp 1668240031
transform 1 0 15640 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_162
timestamp 1668240031
transform 1 0 16008 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_166
timestamp 1668240031
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_169
timestamp 1668240031
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_191
timestamp 1668240031
transform 1 0 18676 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_204
timestamp 1668240031
transform 1 0 19872 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_208
timestamp 1668240031
transform 1 0 20240 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_218
timestamp 1668240031
transform 1 0 21160 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_225
timestamp 1668240031
transform 1 0 21804 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_247
timestamp 1668240031
transform 1 0 23828 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_254
timestamp 1668240031
transform 1 0 24472 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_267
timestamp 1668240031
transform 1 0 25668 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_274
timestamp 1668240031
transform 1 0 26312 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_281
timestamp 1668240031
transform 1 0 26956 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_289
timestamp 1668240031
transform 1 0 27692 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_297
timestamp 1668240031
transform 1 0 28428 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_306
timestamp 1668240031
transform 1 0 29256 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_334
timestamp 1668240031
transform 1 0 31832 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_337
timestamp 1668240031
transform 1 0 32108 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_343
timestamp 1668240031
transform 1 0 32660 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_350
timestamp 1668240031
transform 1 0 33304 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_354
timestamp 1668240031
transform 1 0 33672 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_375
timestamp 1668240031
transform 1 0 35604 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_387
timestamp 1668240031
transform 1 0 36708 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1668240031
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_393
timestamp 1668240031
transform 1 0 37260 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1668240031
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1668240031
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1668240031
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1668240031
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1668240031
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_74
timestamp 1668240031
transform 1 0 7912 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_82
timestamp 1668240031
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_85
timestamp 1668240031
transform 1 0 8924 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_107
timestamp 1668240031
transform 1 0 10948 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_120
timestamp 1668240031
transform 1 0 12144 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_131
timestamp 1668240031
transform 1 0 13156 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_138
timestamp 1668240031
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_141
timestamp 1668240031
transform 1 0 14076 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_146
timestamp 1668240031
transform 1 0 14536 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_159
timestamp 1668240031
transform 1 0 15732 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_169
timestamp 1668240031
transform 1 0 16652 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_182
timestamp 1668240031
transform 1 0 17848 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_190
timestamp 1668240031
transform 1 0 18584 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1668240031
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_197
timestamp 1668240031
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_219
timestamp 1668240031
transform 1 0 21252 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_229
timestamp 1668240031
transform 1 0 22172 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_235
timestamp 1668240031
transform 1 0 22724 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_239
timestamp 1668240031
transform 1 0 23092 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_250
timestamp 1668240031
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1668240031
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_275
timestamp 1668240031
transform 1 0 26404 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_282
timestamp 1668240031
transform 1 0 27048 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_299
timestamp 1668240031
transform 1 0 28612 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_306
timestamp 1668240031
transform 1 0 29256 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_309
timestamp 1668240031
transform 1 0 29532 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_315
timestamp 1668240031
transform 1 0 30084 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_326
timestamp 1668240031
transform 1 0 31096 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_340
timestamp 1668240031
transform 1 0 32384 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_347
timestamp 1668240031
transform 1 0 33028 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_359
timestamp 1668240031
transform 1 0 34132 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1668240031
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_365
timestamp 1668240031
transform 1 0 34684 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_370
timestamp 1668240031
transform 1 0 35144 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_382
timestamp 1668240031
transform 1 0 36248 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1668240031
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1668240031
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1668240031
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1668240031
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1668240031
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1668240031
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1668240031
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_69
timestamp 1668240031
transform 1 0 7452 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_95
timestamp 1668240031
transform 1 0 9844 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_108
timestamp 1668240031
transform 1 0 11040 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_113
timestamp 1668240031
transform 1 0 11500 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_118
timestamp 1668240031
transform 1 0 11960 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_125
timestamp 1668240031
transform 1 0 12604 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_138
timestamp 1668240031
transform 1 0 13800 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_166
timestamp 1668240031
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_169
timestamp 1668240031
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_180
timestamp 1668240031
transform 1 0 17664 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_184
timestamp 1668240031
transform 1 0 18032 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_205
timestamp 1668240031
transform 1 0 19964 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_211
timestamp 1668240031
transform 1 0 20516 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_221
timestamp 1668240031
transform 1 0 21436 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_225
timestamp 1668240031
transform 1 0 21804 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_248
timestamp 1668240031
transform 1 0 23920 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_254
timestamp 1668240031
transform 1 0 24472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_264
timestamp 1668240031
transform 1 0 25392 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_31_277
timestamp 1668240031
transform 1 0 26588 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_281
timestamp 1668240031
transform 1 0 26956 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_303
timestamp 1668240031
transform 1 0 28980 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_310
timestamp 1668240031
transform 1 0 29624 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_325
timestamp 1668240031
transform 1 0 31004 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_333
timestamp 1668240031
transform 1 0 31740 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_337
timestamp 1668240031
transform 1 0 32108 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_359
timestamp 1668240031
transform 1 0 34132 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_371
timestamp 1668240031
transform 1 0 35236 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_383
timestamp 1668240031
transform 1 0 36340 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1668240031
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_393
timestamp 1668240031
transform 1 0 37260 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1668240031
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1668240031
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1668240031
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1668240031
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1668240031
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1668240031
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1668240031
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_77
timestamp 1668240031
transform 1 0 8188 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_82
timestamp 1668240031
transform 1 0 8648 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_85
timestamp 1668240031
transform 1 0 8924 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_90
timestamp 1668240031
transform 1 0 9384 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_94
timestamp 1668240031
transform 1 0 9752 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_104
timestamp 1668240031
transform 1 0 10672 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_117
timestamp 1668240031
transform 1 0 11868 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_121
timestamp 1668240031
transform 1 0 12236 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_125
timestamp 1668240031
transform 1 0 12604 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_138
timestamp 1668240031
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_141
timestamp 1668240031
transform 1 0 14076 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_152
timestamp 1668240031
transform 1 0 15088 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_161
timestamp 1668240031
transform 1 0 15916 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_185
timestamp 1668240031
transform 1 0 18124 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1668240031
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_197
timestamp 1668240031
transform 1 0 19228 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_202
timestamp 1668240031
transform 1 0 19688 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_32_230
timestamp 1668240031
transform 1 0 22264 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_238
timestamp 1668240031
transform 1 0 23000 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_250
timestamp 1668240031
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_253
timestamp 1668240031
transform 1 0 24380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_258
timestamp 1668240031
transform 1 0 24840 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_264
timestamp 1668240031
transform 1 0 25392 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_274
timestamp 1668240031
transform 1 0 26312 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_298
timestamp 1668240031
transform 1 0 28520 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_306
timestamp 1668240031
transform 1 0 29256 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_309
timestamp 1668240031
transform 1 0 29532 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_332
timestamp 1668240031
transform 1 0 31648 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_340
timestamp 1668240031
transform 1 0 32384 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_362
timestamp 1668240031
transform 1 0 34408 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1668240031
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_377
timestamp 1668240031
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_389
timestamp 1668240031
transform 1 0 36892 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_393
timestamp 1668240031
transform 1 0 37260 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1668240031
transform 1 0 1380 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_8
timestamp 1668240031
transform 1 0 1840 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_20
timestamp 1668240031
transform 1 0 2944 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_32
timestamp 1668240031
transform 1 0 4048 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_44
timestamp 1668240031
transform 1 0 5152 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_57
timestamp 1668240031
transform 1 0 6348 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_65
timestamp 1668240031
transform 1 0 7084 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_71
timestamp 1668240031
transform 1 0 7636 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_84
timestamp 1668240031
transform 1 0 8832 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1668240031
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_113
timestamp 1668240031
transform 1 0 11500 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_135
timestamp 1668240031
transform 1 0 13524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1668240031
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1668240031
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_169
timestamp 1668240031
transform 1 0 16652 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_174
timestamp 1668240031
transform 1 0 17112 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_181
timestamp 1668240031
transform 1 0 17756 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_189
timestamp 1668240031
transform 1 0 18492 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_193
timestamp 1668240031
transform 1 0 18860 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_206
timestamp 1668240031
transform 1 0 20056 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_215
timestamp 1668240031
transform 1 0 20884 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_222
timestamp 1668240031
transform 1 0 21528 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_225
timestamp 1668240031
transform 1 0 21804 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_234
timestamp 1668240031
transform 1 0 22632 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_258
timestamp 1668240031
transform 1 0 24840 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_271
timestamp 1668240031
transform 1 0 26036 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_278
timestamp 1668240031
transform 1 0 26680 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_281
timestamp 1668240031
transform 1 0 26956 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_292
timestamp 1668240031
transform 1 0 27968 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_299
timestamp 1668240031
transform 1 0 28612 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_307
timestamp 1668240031
transform 1 0 29348 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_317
timestamp 1668240031
transform 1 0 30268 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_324
timestamp 1668240031
transform 1 0 30912 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_331
timestamp 1668240031
transform 1 0 31556 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1668240031
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_337
timestamp 1668240031
transform 1 0 32108 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_342
timestamp 1668240031
transform 1 0 32568 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_357
timestamp 1668240031
transform 1 0 33948 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_364
timestamp 1668240031
transform 1 0 34592 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_371
timestamp 1668240031
transform 1 0 35236 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_378
timestamp 1668240031
transform 1 0 35880 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_386
timestamp 1668240031
transform 1 0 36616 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_390
timestamp 1668240031
transform 1 0 36984 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_393
timestamp 1668240031
transform 1 0 37260 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1668240031
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1668240031
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1668240031
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1668240031
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1668240031
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_53
timestamp 1668240031
transform 1 0 5980 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_61
timestamp 1668240031
transform 1 0 6716 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_82
timestamp 1668240031
transform 1 0 8648 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_85
timestamp 1668240031
transform 1 0 8924 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_96
timestamp 1668240031
transform 1 0 9936 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_104
timestamp 1668240031
transform 1 0 10672 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_108
timestamp 1668240031
transform 1 0 11040 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_115
timestamp 1668240031
transform 1 0 11684 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_128
timestamp 1668240031
transform 1 0 12880 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_141
timestamp 1668240031
transform 1 0 14076 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_146
timestamp 1668240031
transform 1 0 14536 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_152
timestamp 1668240031
transform 1 0 15088 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_156
timestamp 1668240031
transform 1 0 15456 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_160
timestamp 1668240031
transform 1 0 15824 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_181
timestamp 1668240031
transform 1 0 17756 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_187
timestamp 1668240031
transform 1 0 18308 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_194
timestamp 1668240031
transform 1 0 18952 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_197
timestamp 1668240031
transform 1 0 19228 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_221
timestamp 1668240031
transform 1 0 21436 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_234
timestamp 1668240031
transform 1 0 22632 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_244
timestamp 1668240031
transform 1 0 23552 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_253
timestamp 1668240031
transform 1 0 24380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_264
timestamp 1668240031
transform 1 0 25392 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_277
timestamp 1668240031
transform 1 0 26588 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_283
timestamp 1668240031
transform 1 0 27140 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_290
timestamp 1668240031
transform 1 0 27784 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_298
timestamp 1668240031
transform 1 0 28520 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_306
timestamp 1668240031
transform 1 0 29256 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_309
timestamp 1668240031
transform 1 0 29532 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_315
timestamp 1668240031
transform 1 0 30084 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_337
timestamp 1668240031
transform 1 0 32108 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_347
timestamp 1668240031
transform 1 0 33028 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_360
timestamp 1668240031
transform 1 0 34224 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_365
timestamp 1668240031
transform 1 0 34684 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_376
timestamp 1668240031
transform 1 0 35696 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_388
timestamp 1668240031
transform 1 0 36800 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1668240031
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1668240031
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_27
timestamp 1668240031
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_39
timestamp 1668240031
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1668240031
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1668240031
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1668240031
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_69
timestamp 1668240031
transform 1 0 7452 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_76
timestamp 1668240031
transform 1 0 8096 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_88
timestamp 1668240031
transform 1 0 9200 0 -1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_35_99
timestamp 1668240031
transform 1 0 10212 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1668240031
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_113
timestamp 1668240031
transform 1 0 11500 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_117
timestamp 1668240031
transform 1 0 11868 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_121
timestamp 1668240031
transform 1 0 12236 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_129
timestamp 1668240031
transform 1 0 12972 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_140
timestamp 1668240031
transform 1 0 13984 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_146
timestamp 1668240031
transform 1 0 14536 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_150
timestamp 1668240031
transform 1 0 14904 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_158
timestamp 1668240031
transform 1 0 15640 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_166
timestamp 1668240031
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_169
timestamp 1668240031
transform 1 0 16652 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_175
timestamp 1668240031
transform 1 0 17204 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_182
timestamp 1668240031
transform 1 0 17848 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_206
timestamp 1668240031
transform 1 0 20056 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_219
timestamp 1668240031
transform 1 0 21252 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1668240031
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_225
timestamp 1668240031
transform 1 0 21804 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_236
timestamp 1668240031
transform 1 0 22816 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_247
timestamp 1668240031
transform 1 0 23828 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_254
timestamp 1668240031
transform 1 0 24472 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_271
timestamp 1668240031
transform 1 0 26036 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_278
timestamp 1668240031
transform 1 0 26680 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_281
timestamp 1668240031
transform 1 0 26956 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_303
timestamp 1668240031
transform 1 0 28980 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_311
timestamp 1668240031
transform 1 0 29716 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_324
timestamp 1668240031
transform 1 0 30912 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_337
timestamp 1668240031
transform 1 0 32108 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_346
timestamp 1668240031
transform 1 0 32936 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_352
timestamp 1668240031
transform 1 0 33488 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_360
timestamp 1668240031
transform 1 0 34224 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_389
timestamp 1668240031
transform 1 0 36892 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_35_393
timestamp 1668240031
transform 1 0 37260 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1668240031
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1668240031
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1668240031
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1668240031
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1668240031
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1668240031
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_65
timestamp 1668240031
transform 1 0 7084 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_70
timestamp 1668240031
transform 1 0 7544 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1668240031
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1668240031
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_85
timestamp 1668240031
transform 1 0 8924 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_92
timestamp 1668240031
transform 1 0 9568 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_99
timestamp 1668240031
transform 1 0 10212 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_106
timestamp 1668240031
transform 1 0 10856 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_114
timestamp 1668240031
transform 1 0 11592 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_120
timestamp 1668240031
transform 1 0 12144 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1668240031
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1668240031
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_141
timestamp 1668240031
transform 1 0 14076 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_163
timestamp 1668240031
transform 1 0 16100 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_167
timestamp 1668240031
transform 1 0 16468 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_171
timestamp 1668240031
transform 1 0 16836 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_181
timestamp 1668240031
transform 1 0 17756 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_194
timestamp 1668240031
transform 1 0 18952 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_197
timestamp 1668240031
transform 1 0 19228 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_201
timestamp 1668240031
transform 1 0 19596 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_205
timestamp 1668240031
transform 1 0 19964 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_229
timestamp 1668240031
transform 1 0 22172 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_237
timestamp 1668240031
transform 1 0 22908 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_243
timestamp 1668240031
transform 1 0 23460 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_250
timestamp 1668240031
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_253
timestamp 1668240031
transform 1 0 24380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_258
timestamp 1668240031
transform 1 0 24840 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_275
timestamp 1668240031
transform 1 0 26404 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_279
timestamp 1668240031
transform 1 0 26772 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_283
timestamp 1668240031
transform 1 0 27140 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_290
timestamp 1668240031
transform 1 0 27784 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_298
timestamp 1668240031
transform 1 0 28520 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_306
timestamp 1668240031
transform 1 0 29256 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_309
timestamp 1668240031
transform 1 0 29532 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_318
timestamp 1668240031
transform 1 0 30360 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_324
timestamp 1668240031
transform 1 0 30912 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_330
timestamp 1668240031
transform 1 0 31464 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_341
timestamp 1668240031
transform 1 0 32476 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_349
timestamp 1668240031
transform 1 0 33212 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_358
timestamp 1668240031
transform 1 0 34040 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_36_365
timestamp 1668240031
transform 1 0 34684 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_372
timestamp 1668240031
transform 1 0 35328 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_378
timestamp 1668240031
transform 1 0 35880 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_382
timestamp 1668240031
transform 1 0 36248 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_386
timestamp 1668240031
transform 1 0 36616 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_390
timestamp 1668240031
transform 1 0 36984 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1668240031
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1668240031
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_27
timestamp 1668240031
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_39
timestamp 1668240031
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1668240031
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1668240031
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_37_57
timestamp 1668240031
transform 1 0 6348 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_37_80
timestamp 1668240031
transform 1 0 8464 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_86
timestamp 1668240031
transform 1 0 9016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_107
timestamp 1668240031
transform 1 0 10948 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1668240031
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_113
timestamp 1668240031
transform 1 0 11500 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_135
timestamp 1668240031
transform 1 0 13524 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_142
timestamp 1668240031
transform 1 0 14168 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_148
timestamp 1668240031
transform 1 0 14720 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_155
timestamp 1668240031
transform 1 0 15364 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_166
timestamp 1668240031
transform 1 0 16376 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_169
timestamp 1668240031
transform 1 0 16652 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_191
timestamp 1668240031
transform 1 0 18676 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_195
timestamp 1668240031
transform 1 0 19044 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_199
timestamp 1668240031
transform 1 0 19412 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_37_216
timestamp 1668240031
transform 1 0 20976 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_225
timestamp 1668240031
transform 1 0 21804 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_230
timestamp 1668240031
transform 1 0 22264 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_234
timestamp 1668240031
transform 1 0 22632 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_255
timestamp 1668240031
transform 1 0 24564 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_268
timestamp 1668240031
transform 1 0 25760 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_275
timestamp 1668240031
transform 1 0 26404 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1668240031
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_281
timestamp 1668240031
transform 1 0 26956 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_303
timestamp 1668240031
transform 1 0 28980 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_316
timestamp 1668240031
transform 1 0 30176 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_323
timestamp 1668240031
transform 1 0 30820 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1668240031
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_337
timestamp 1668240031
transform 1 0 32108 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_347
timestamp 1668240031
transform 1 0 33028 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_351
timestamp 1668240031
transform 1 0 33396 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_372
timestamp 1668240031
transform 1 0 35328 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_379
timestamp 1668240031
transform 1 0 35972 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_386
timestamp 1668240031
transform 1 0 36616 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_393
timestamp 1668240031
transform 1 0 37260 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1668240031
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1668240031
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1668240031
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1668240031
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1668240031
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_56
timestamp 1668240031
transform 1 0 6256 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_69
timestamp 1668240031
transform 1 0 7452 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_82
timestamp 1668240031
transform 1 0 8648 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_85
timestamp 1668240031
transform 1 0 8924 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_96
timestamp 1668240031
transform 1 0 9936 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_122
timestamp 1668240031
transform 1 0 12328 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_135
timestamp 1668240031
transform 1 0 13524 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1668240031
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_38_141
timestamp 1668240031
transform 1 0 14076 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_164
timestamp 1668240031
transform 1 0 16192 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_171
timestamp 1668240031
transform 1 0 16836 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_178
timestamp 1668240031
transform 1 0 17480 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_186
timestamp 1668240031
transform 1 0 18216 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_192
timestamp 1668240031
transform 1 0 18768 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_38_197
timestamp 1668240031
transform 1 0 19228 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_38_209
timestamp 1668240031
transform 1 0 20332 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_215
timestamp 1668240031
transform 1 0 20884 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_225
timestamp 1668240031
transform 1 0 21804 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_229
timestamp 1668240031
transform 1 0 22172 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_250
timestamp 1668240031
transform 1 0 24104 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_253
timestamp 1668240031
transform 1 0 24380 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_259
timestamp 1668240031
transform 1 0 24932 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_269
timestamp 1668240031
transform 1 0 25852 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_273
timestamp 1668240031
transform 1 0 26220 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_277
timestamp 1668240031
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_292
timestamp 1668240031
transform 1 0 27968 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_296
timestamp 1668240031
transform 1 0 28336 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_304
timestamp 1668240031
transform 1 0 29072 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_309
timestamp 1668240031
transform 1 0 29532 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_314
timestamp 1668240031
transform 1 0 29992 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_321
timestamp 1668240031
transform 1 0 30636 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_347
timestamp 1668240031
transform 1 0 33028 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_356
timestamp 1668240031
transform 1 0 33856 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_365
timestamp 1668240031
transform 1 0 34684 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_390
timestamp 1668240031
transform 1 0 36984 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1668240031
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1668240031
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1668240031
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1668240031
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1668240031
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1668240031
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_57
timestamp 1668240031
transform 1 0 6348 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_63
timestamp 1668240031
transform 1 0 6900 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_84
timestamp 1668240031
transform 1 0 8832 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_97
timestamp 1668240031
transform 1 0 10028 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_110
timestamp 1668240031
transform 1 0 11224 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_113
timestamp 1668240031
transform 1 0 11500 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_125
timestamp 1668240031
transform 1 0 12604 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_149
timestamp 1668240031
transform 1 0 14812 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1668240031
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1668240031
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_169
timestamp 1668240031
transform 1 0 16652 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_174
timestamp 1668240031
transform 1 0 17112 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_198
timestamp 1668240031
transform 1 0 19320 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_222
timestamp 1668240031
transform 1 0 21528 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_225
timestamp 1668240031
transform 1 0 21804 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_233
timestamp 1668240031
transform 1 0 22540 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_241
timestamp 1668240031
transform 1 0 23276 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_39_258
timestamp 1668240031
transform 1 0 24840 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_266
timestamp 1668240031
transform 1 0 25576 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_277
timestamp 1668240031
transform 1 0 26588 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_281
timestamp 1668240031
transform 1 0 26956 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_303
timestamp 1668240031
transform 1 0 28980 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_332
timestamp 1668240031
transform 1 0 31648 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_337
timestamp 1668240031
transform 1 0 32108 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_346
timestamp 1668240031
transform 1 0 32936 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_357
timestamp 1668240031
transform 1 0 33948 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_361
timestamp 1668240031
transform 1 0 34316 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_365
timestamp 1668240031
transform 1 0 34684 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_390
timestamp 1668240031
transform 1 0 36984 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_393
timestamp 1668240031
transform 1 0 37260 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_3
timestamp 1668240031
transform 1 0 1380 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_8
timestamp 1668240031
transform 1 0 1840 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_20
timestamp 1668240031
transform 1 0 2944 0 1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1668240031
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1668240031
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1668240031
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_65
timestamp 1668240031
transform 1 0 7084 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_69
timestamp 1668240031
transform 1 0 7452 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_82
timestamp 1668240031
transform 1 0 8648 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_85
timestamp 1668240031
transform 1 0 8924 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_93
timestamp 1668240031
transform 1 0 9660 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_107
timestamp 1668240031
transform 1 0 10948 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_114
timestamp 1668240031
transform 1 0 11592 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_129
timestamp 1668240031
transform 1 0 12972 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_136
timestamp 1668240031
transform 1 0 13616 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_141
timestamp 1668240031
transform 1 0 14076 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_146
timestamp 1668240031
transform 1 0 14536 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_150
timestamp 1668240031
transform 1 0 14904 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_154
timestamp 1668240031
transform 1 0 15272 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_178
timestamp 1668240031
transform 1 0 17480 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_184
timestamp 1668240031
transform 1 0 18032 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_188
timestamp 1668240031
transform 1 0 18400 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_197
timestamp 1668240031
transform 1 0 19228 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_210
timestamp 1668240031
transform 1 0 20424 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_216
timestamp 1668240031
transform 1 0 20976 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_220
timestamp 1668240031
transform 1 0 21344 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_232
timestamp 1668240031
transform 1 0 22448 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_236
timestamp 1668240031
transform 1 0 22816 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_240
timestamp 1668240031
transform 1 0 23184 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_247
timestamp 1668240031
transform 1 0 23828 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1668240031
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_253
timestamp 1668240031
transform 1 0 24380 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_270
timestamp 1668240031
transform 1 0 25944 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_283
timestamp 1668240031
transform 1 0 27140 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_295
timestamp 1668240031
transform 1 0 28244 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_306
timestamp 1668240031
transform 1 0 29256 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_309
timestamp 1668240031
transform 1 0 29532 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_334
timestamp 1668240031
transform 1 0 31832 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_345
timestamp 1668240031
transform 1 0 32844 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_351
timestamp 1668240031
transform 1 0 33396 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_360
timestamp 1668240031
transform 1 0 34224 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_365
timestamp 1668240031
transform 1 0 34684 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_376
timestamp 1668240031
transform 1 0 35696 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_388
timestamp 1668240031
transform 1 0 36800 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_392
timestamp 1668240031
transform 1 0 37168 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1668240031
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1668240031
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_27
timestamp 1668240031
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_39
timestamp 1668240031
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1668240031
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1668240031
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1668240031
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_89
timestamp 1668240031
transform 1 0 9292 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_93
timestamp 1668240031
transform 1 0 9660 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_97
timestamp 1668240031
transform 1 0 10028 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_110
timestamp 1668240031
transform 1 0 11224 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_113
timestamp 1668240031
transform 1 0 11500 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_124
timestamp 1668240031
transform 1 0 12512 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_137
timestamp 1668240031
transform 1 0 13708 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_145
timestamp 1668240031
transform 1 0 14444 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_151
timestamp 1668240031
transform 1 0 14996 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_158
timestamp 1668240031
transform 1 0 15640 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_162
timestamp 1668240031
transform 1 0 16008 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_166
timestamp 1668240031
transform 1 0 16376 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_169
timestamp 1668240031
transform 1 0 16652 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_177
timestamp 1668240031
transform 1 0 17388 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_184
timestamp 1668240031
transform 1 0 18032 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_190
timestamp 1668240031
transform 1 0 18584 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_200
timestamp 1668240031
transform 1 0 19504 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_204
timestamp 1668240031
transform 1 0 19872 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_208
timestamp 1668240031
transform 1 0 20240 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_41_221
timestamp 1668240031
transform 1 0 21436 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_225
timestamp 1668240031
transform 1 0 21804 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_247
timestamp 1668240031
transform 1 0 23828 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_271
timestamp 1668240031
transform 1 0 26036 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_278
timestamp 1668240031
transform 1 0 26680 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_281
timestamp 1668240031
transform 1 0 26956 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_286
timestamp 1668240031
transform 1 0 27416 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_293
timestamp 1668240031
transform 1 0 28060 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_299
timestamp 1668240031
transform 1 0 28612 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_307
timestamp 1668240031
transform 1 0 29348 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_316
timestamp 1668240031
transform 1 0 30176 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_323
timestamp 1668240031
transform 1 0 30820 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_330
timestamp 1668240031
transform 1 0 31464 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_41_337
timestamp 1668240031
transform 1 0 32108 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_343
timestamp 1668240031
transform 1 0 32660 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_349
timestamp 1668240031
transform 1 0 33212 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_358
timestamp 1668240031
transform 1 0 34040 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_371
timestamp 1668240031
transform 1 0 35236 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_386
timestamp 1668240031
transform 1 0 36616 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_393
timestamp 1668240031
transform 1 0 37260 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1668240031
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1668240031
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1668240031
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1668240031
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1668240031
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1668240031
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_65
timestamp 1668240031
transform 1 0 7084 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_71
timestamp 1668240031
transform 1 0 7636 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_75
timestamp 1668240031
transform 1 0 8004 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_82
timestamp 1668240031
transform 1 0 8648 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_85
timestamp 1668240031
transform 1 0 8924 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_98
timestamp 1668240031
transform 1 0 10120 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_105
timestamp 1668240031
transform 1 0 10764 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_129
timestamp 1668240031
transform 1 0 12972 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_137
timestamp 1668240031
transform 1 0 13708 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_42_141
timestamp 1668240031
transform 1 0 14076 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_163
timestamp 1668240031
transform 1 0 16100 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_167
timestamp 1668240031
transform 1 0 16468 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_188
timestamp 1668240031
transform 1 0 18400 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_197
timestamp 1668240031
transform 1 0 19228 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_208
timestamp 1668240031
transform 1 0 20240 0 1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_42_217
timestamp 1668240031
transform 1 0 21068 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_229
timestamp 1668240031
transform 1 0 22172 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_42_235
timestamp 1668240031
transform 1 0 22724 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_42_250
timestamp 1668240031
transform 1 0 24104 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_253
timestamp 1668240031
transform 1 0 24380 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_264
timestamp 1668240031
transform 1 0 25392 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_271
timestamp 1668240031
transform 1 0 26036 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_42_297
timestamp 1668240031
transform 1 0 28428 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_305
timestamp 1668240031
transform 1 0 29164 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_42_309
timestamp 1668240031
transform 1 0 29532 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_325
timestamp 1668240031
transform 1 0 31004 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_334
timestamp 1668240031
transform 1 0 31832 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_343
timestamp 1668240031
transform 1 0 32660 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_354
timestamp 1668240031
transform 1 0 33672 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_42_361
timestamp 1668240031
transform 1 0 34316 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_42_365
timestamp 1668240031
transform 1 0 34684 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_372
timestamp 1668240031
transform 1 0 35328 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_379
timestamp 1668240031
transform 1 0 35972 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_386
timestamp 1668240031
transform 1 0 36616 0 1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1668240031
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1668240031
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1668240031
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1668240031
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1668240031
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1668240031
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1668240031
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_69
timestamp 1668240031
transform 1 0 7452 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_77
timestamp 1668240031
transform 1 0 8188 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_43_82
timestamp 1668240031
transform 1 0 8648 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_108
timestamp 1668240031
transform 1 0 11040 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_113
timestamp 1668240031
transform 1 0 11500 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_119
timestamp 1668240031
transform 1 0 12052 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_123
timestamp 1668240031
transform 1 0 12420 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_131
timestamp 1668240031
transform 1 0 13156 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_135
timestamp 1668240031
transform 1 0 13524 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_159
timestamp 1668240031
transform 1 0 15732 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_166
timestamp 1668240031
transform 1 0 16376 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_169
timestamp 1668240031
transform 1 0 16652 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_191
timestamp 1668240031
transform 1 0 18676 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_198
timestamp 1668240031
transform 1 0 19320 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_222
timestamp 1668240031
transform 1 0 21528 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_43_225
timestamp 1668240031
transform 1 0 21804 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_43_248
timestamp 1668240031
transform 1 0 23920 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_263
timestamp 1668240031
transform 1 0 25300 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_276
timestamp 1668240031
transform 1 0 26496 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_281
timestamp 1668240031
transform 1 0 26956 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_303
timestamp 1668240031
transform 1 0 28980 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_314
timestamp 1668240031
transform 1 0 29992 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_322
timestamp 1668240031
transform 1 0 30728 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 1668240031
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1668240031
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_337
timestamp 1668240031
transform 1 0 32108 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_345
timestamp 1668240031
transform 1 0 32844 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_349
timestamp 1668240031
transform 1 0 33212 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_356
timestamp 1668240031
transform 1 0 33856 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1668240031
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1668240031
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_43_393
timestamp 1668240031
transform 1 0 37260 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1668240031
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1668240031
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1668240031
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1668240031
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1668240031
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1668240031
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_65
timestamp 1668240031
transform 1 0 7084 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_71
timestamp 1668240031
transform 1 0 7636 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_75
timestamp 1668240031
transform 1 0 8004 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_82
timestamp 1668240031
transform 1 0 8648 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_85
timestamp 1668240031
transform 1 0 8924 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_44_102
timestamp 1668240031
transform 1 0 10488 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_108
timestamp 1668240031
transform 1 0 11040 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_112
timestamp 1668240031
transform 1 0 11408 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_136
timestamp 1668240031
transform 1 0 13616 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_141
timestamp 1668240031
transform 1 0 14076 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_154
timestamp 1668240031
transform 1 0 15272 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_162
timestamp 1668240031
transform 1 0 16008 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_166
timestamp 1668240031
transform 1 0 16376 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_179
timestamp 1668240031
transform 1 0 17572 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_44_194
timestamp 1668240031
transform 1 0 18952 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_44_197
timestamp 1668240031
transform 1 0 19228 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_209
timestamp 1668240031
transform 1 0 20332 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_233
timestamp 1668240031
transform 1 0 22540 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_239
timestamp 1668240031
transform 1 0 23092 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_44_249
timestamp 1668240031
transform 1 0 24012 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_253
timestamp 1668240031
transform 1 0 24380 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_258
timestamp 1668240031
transform 1 0 24840 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_265
timestamp 1668240031
transform 1 0 25484 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_278
timestamp 1668240031
transform 1 0 26680 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_285
timestamp 1668240031
transform 1 0 27324 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_292
timestamp 1668240031
transform 1 0 27968 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_303
timestamp 1668240031
transform 1 0 28980 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1668240031
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_309
timestamp 1668240031
transform 1 0 29532 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_44_336
timestamp 1668240031
transform 1 0 32016 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_342
timestamp 1668240031
transform 1 0 32568 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_351
timestamp 1668240031
transform 1 0 33396 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_362
timestamp 1668240031
transform 1 0 34408 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_365
timestamp 1668240031
transform 1 0 34684 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_44_392
timestamp 1668240031
transform 1 0 37168 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1668240031
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1668240031
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1668240031
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1668240031
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1668240031
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1668240031
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_57
timestamp 1668240031
transform 1 0 6348 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_65
timestamp 1668240031
transform 1 0 7084 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_88
timestamp 1668240031
transform 1 0 9200 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_101
timestamp 1668240031
transform 1 0 10396 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_45_110
timestamp 1668240031
transform 1 0 11224 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_113
timestamp 1668240031
transform 1 0 11500 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_45_124
timestamp 1668240031
transform 1 0 12512 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_152
timestamp 1668240031
transform 1 0 15088 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_45_165
timestamp 1668240031
transform 1 0 16284 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_169
timestamp 1668240031
transform 1 0 16652 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_176
timestamp 1668240031
transform 1 0 17296 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_182
timestamp 1668240031
transform 1 0 17848 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_203
timestamp 1668240031
transform 1 0 19780 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_207
timestamp 1668240031
transform 1 0 20148 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_219
timestamp 1668240031
transform 1 0 21252 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1668240031
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_225
timestamp 1668240031
transform 1 0 21804 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_45_230
timestamp 1668240031
transform 1 0 22264 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_45_247
timestamp 1668240031
transform 1 0 23828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_262
timestamp 1668240031
transform 1 0 25208 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_269
timestamp 1668240031
transform 1 0 25852 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_276
timestamp 1668240031
transform 1 0 26496 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_281
timestamp 1668240031
transform 1 0 26956 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_45_289
timestamp 1668240031
transform 1 0 27692 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_295
timestamp 1668240031
transform 1 0 28244 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_301
timestamp 1668240031
transform 1 0 28796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_308
timestamp 1668240031
transform 1 0 29440 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_316
timestamp 1668240031
transform 1 0 30176 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_327
timestamp 1668240031
transform 1 0 31188 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_334
timestamp 1668240031
transform 1 0 31832 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_337
timestamp 1668240031
transform 1 0 32108 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_346
timestamp 1668240031
transform 1 0 32936 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_353
timestamp 1668240031
transform 1 0 33580 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_359
timestamp 1668240031
transform 1 0 34132 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_369
timestamp 1668240031
transform 1 0 35052 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_380
timestamp 1668240031
transform 1 0 36064 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_387
timestamp 1668240031
transform 1 0 36708 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1668240031
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_45_393
timestamp 1668240031
transform 1 0 37260 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1668240031
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1668240031
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1668240031
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1668240031
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1668240031
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1668240031
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_65
timestamp 1668240031
transform 1 0 7084 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_69
timestamp 1668240031
transform 1 0 7452 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_82
timestamp 1668240031
transform 1 0 8648 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_85
timestamp 1668240031
transform 1 0 8924 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_91
timestamp 1668240031
transform 1 0 9476 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_95
timestamp 1668240031
transform 1 0 9844 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_122
timestamp 1668240031
transform 1 0 12328 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_135
timestamp 1668240031
transform 1 0 13524 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1668240031
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_46_141
timestamp 1668240031
transform 1 0 14076 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_46_147
timestamp 1668240031
transform 1 0 14628 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_156
timestamp 1668240031
transform 1 0 15456 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_180
timestamp 1668240031
transform 1 0 17664 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_184
timestamp 1668240031
transform 1 0 18032 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_194
timestamp 1668240031
transform 1 0 18952 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_197
timestamp 1668240031
transform 1 0 19228 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_208
timestamp 1668240031
transform 1 0 20240 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_215
timestamp 1668240031
transform 1 0 20884 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_222
timestamp 1668240031
transform 1 0 21528 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_228
timestamp 1668240031
transform 1 0 22080 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_238
timestamp 1668240031
transform 1 0 23000 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1668240031
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1668240031
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_253
timestamp 1668240031
transform 1 0 24380 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_279
timestamp 1668240031
transform 1 0 26772 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_303
timestamp 1668240031
transform 1 0 28980 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1668240031
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_309
timestamp 1668240031
transform 1 0 29532 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_315
timestamp 1668240031
transform 1 0 30084 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_323
timestamp 1668240031
transform 1 0 30820 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_332
timestamp 1668240031
transform 1 0 31648 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_345
timestamp 1668240031
transform 1 0 32844 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_349
timestamp 1668240031
transform 1 0 33212 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1668240031
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1668240031
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_365
timestamp 1668240031
transform 1 0 34684 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_376
timestamp 1668240031
transform 1 0 35696 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_383
timestamp 1668240031
transform 1 0 36340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_46_392
timestamp 1668240031
transform 1 0 37168 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_3
timestamp 1668240031
transform 1 0 1380 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_8
timestamp 1668240031
transform 1 0 1840 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_20
timestamp 1668240031
transform 1 0 2944 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_32
timestamp 1668240031
transform 1 0 4048 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_44
timestamp 1668240031
transform 1 0 5152 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_57
timestamp 1668240031
transform 1 0 6348 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_79
timestamp 1668240031
transform 1 0 8372 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_86
timestamp 1668240031
transform 1 0 9016 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_110
timestamp 1668240031
transform 1 0 11224 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_113
timestamp 1668240031
transform 1 0 11500 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_118
timestamp 1668240031
transform 1 0 11960 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_131
timestamp 1668240031
transform 1 0 13156 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_138
timestamp 1668240031
transform 1 0 13800 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_151
timestamp 1668240031
transform 1 0 14996 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_164
timestamp 1668240031
transform 1 0 16192 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_169
timestamp 1668240031
transform 1 0 16652 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_180
timestamp 1668240031
transform 1 0 17664 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_187
timestamp 1668240031
transform 1 0 18308 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_211
timestamp 1668240031
transform 1 0 20516 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_218
timestamp 1668240031
transform 1 0 21160 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_47_225
timestamp 1668240031
transform 1 0 21804 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_47_230
timestamp 1668240031
transform 1 0 22264 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_236
timestamp 1668240031
transform 1 0 22816 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_243
timestamp 1668240031
transform 1 0 23460 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_256
timestamp 1668240031
transform 1 0 24656 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_269
timestamp 1668240031
transform 1 0 25852 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_47_278
timestamp 1668240031
transform 1 0 26680 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_281
timestamp 1668240031
transform 1 0 26956 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_47_296
timestamp 1668240031
transform 1 0 28336 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_307
timestamp 1668240031
transform 1 0 29348 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_317
timestamp 1668240031
transform 1 0 30268 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_328
timestamp 1668240031
transform 1 0 31280 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_337
timestamp 1668240031
transform 1 0 32108 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_345
timestamp 1668240031
transform 1 0 32844 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_349
timestamp 1668240031
transform 1 0 33212 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_353
timestamp 1668240031
transform 1 0 33580 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_360
timestamp 1668240031
transform 1 0 34224 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_366
timestamp 1668240031
transform 1 0 34776 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_388
timestamp 1668240031
transform 1 0 36800 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_393
timestamp 1668240031
transform 1 0 37260 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1668240031
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1668240031
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1668240031
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1668240031
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1668240031
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_53
timestamp 1668240031
transform 1 0 5980 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_61
timestamp 1668240031
transform 1 0 6716 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_67
timestamp 1668240031
transform 1 0 7268 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_71
timestamp 1668240031
transform 1 0 7636 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_48_81
timestamp 1668240031
transform 1 0 8556 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_48_85
timestamp 1668240031
transform 1 0 8924 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_96
timestamp 1668240031
transform 1 0 9936 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_103
timestamp 1668240031
transform 1 0 10580 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_116
timestamp 1668240031
transform 1 0 11776 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_122
timestamp 1668240031
transform 1 0 12328 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_129
timestamp 1668240031
transform 1 0 12972 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_48_138
timestamp 1668240031
transform 1 0 13800 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_141
timestamp 1668240031
transform 1 0 14076 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_152
timestamp 1668240031
transform 1 0 15088 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_159
timestamp 1668240031
transform 1 0 15732 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_166
timestamp 1668240031
transform 1 0 16376 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_170
timestamp 1668240031
transform 1 0 16744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_180
timestamp 1668240031
transform 1 0 17664 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_184
timestamp 1668240031
transform 1 0 18032 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_194
timestamp 1668240031
transform 1 0 18952 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_197
timestamp 1668240031
transform 1 0 19228 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_206
timestamp 1668240031
transform 1 0 20056 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_230
timestamp 1668240031
transform 1 0 22264 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_238
timestamp 1668240031
transform 1 0 23000 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_48_249
timestamp 1668240031
transform 1 0 24012 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_48_253
timestamp 1668240031
transform 1 0 24380 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_264
timestamp 1668240031
transform 1 0 25392 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_271
timestamp 1668240031
transform 1 0 26036 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_278
timestamp 1668240031
transform 1 0 26680 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_290
timestamp 1668240031
transform 1 0 27784 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_294
timestamp 1668240031
transform 1 0 28152 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_304
timestamp 1668240031
transform 1 0 29072 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_309
timestamp 1668240031
transform 1 0 29532 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_318
timestamp 1668240031
transform 1 0 30360 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_48_342
timestamp 1668240031
transform 1 0 32568 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_48_357
timestamp 1668240031
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1668240031
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_365
timestamp 1668240031
transform 1 0 34684 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_370
timestamp 1668240031
transform 1 0 35144 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_377
timestamp 1668240031
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_389
timestamp 1668240031
transform 1 0 36892 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_393
timestamp 1668240031
transform 1 0 37260 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1668240031
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1668240031
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1668240031
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1668240031
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1668240031
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1668240031
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_57
timestamp 1668240031
transform 1 0 6348 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_79
timestamp 1668240031
transform 1 0 8372 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_87
timestamp 1668240031
transform 1 0 9108 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_49_109
timestamp 1668240031
transform 1 0 11132 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_49_113
timestamp 1668240031
transform 1 0 11500 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_118
timestamp 1668240031
transform 1 0 11960 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_142
timestamp 1668240031
transform 1 0 14168 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_166
timestamp 1668240031
transform 1 0 16376 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_49_169
timestamp 1668240031
transform 1 0 16652 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_195
timestamp 1668240031
transform 1 0 19044 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_202
timestamp 1668240031
transform 1 0 19688 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_209
timestamp 1668240031
transform 1 0 20332 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_217
timestamp 1668240031
transform 1 0 21068 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_222
timestamp 1668240031
transform 1 0 21528 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_49_225
timestamp 1668240031
transform 1 0 21804 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_240
timestamp 1668240031
transform 1 0 23184 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_253
timestamp 1668240031
transform 1 0 24380 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_257
timestamp 1668240031
transform 1 0 24748 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_278
timestamp 1668240031
transform 1 0 26680 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_281
timestamp 1668240031
transform 1 0 26956 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_285
timestamp 1668240031
transform 1 0 27324 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_289
timestamp 1668240031
transform 1 0 27692 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_295
timestamp 1668240031
transform 1 0 28244 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_305
timestamp 1668240031
transform 1 0 29164 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_317
timestamp 1668240031
transform 1 0 30268 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_334
timestamp 1668240031
transform 1 0 31832 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_337
timestamp 1668240031
transform 1 0 32108 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_342
timestamp 1668240031
transform 1 0 32568 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_346
timestamp 1668240031
transform 1 0 32936 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_363
timestamp 1668240031
transform 1 0 34500 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_370
timestamp 1668240031
transform 1 0 35144 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_382
timestamp 1668240031
transform 1 0 36248 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_390
timestamp 1668240031
transform 1 0 36984 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_49_393
timestamp 1668240031
transform 1 0 37260 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1668240031
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1668240031
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1668240031
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1668240031
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_41
timestamp 1668240031
transform 1 0 4876 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_49
timestamp 1668240031
transform 1 0 5612 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_55
timestamp 1668240031
transform 1 0 6164 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_62
timestamp 1668240031
transform 1 0 6808 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_69
timestamp 1668240031
transform 1 0 7452 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_82
timestamp 1668240031
transform 1 0 8648 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_85
timestamp 1668240031
transform 1 0 8924 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_90
timestamp 1668240031
transform 1 0 9384 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_103
timestamp 1668240031
transform 1 0 10580 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_50_129
timestamp 1668240031
transform 1 0 12972 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_50_138
timestamp 1668240031
transform 1 0 13800 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_141
timestamp 1668240031
transform 1 0 14076 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_50_149
timestamp 1668240031
transform 1 0 14812 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_157
timestamp 1668240031
transform 1 0 15548 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_168
timestamp 1668240031
transform 1 0 16560 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_172
timestamp 1668240031
transform 1 0 16928 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_179
timestamp 1668240031
transform 1 0 17572 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_50_194
timestamp 1668240031
transform 1 0 18952 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_197
timestamp 1668240031
transform 1 0 19228 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_50_205
timestamp 1668240031
transform 1 0 19964 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_213
timestamp 1668240031
transform 1 0 20700 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_235
timestamp 1668240031
transform 1 0 22724 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_248
timestamp 1668240031
transform 1 0 23920 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_253
timestamp 1668240031
transform 1 0 24380 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_50_279
timestamp 1668240031
transform 1 0 26772 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_287
timestamp 1668240031
transform 1 0 27508 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_298
timestamp 1668240031
transform 1 0 28520 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_306
timestamp 1668240031
transform 1 0 29256 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_309
timestamp 1668240031
transform 1 0 29532 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_318
timestamp 1668240031
transform 1 0 30360 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_327
timestamp 1668240031
transform 1 0 31188 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_334
timestamp 1668240031
transform 1 0 31832 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_341
timestamp 1668240031
transform 1 0 32476 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_348
timestamp 1668240031
transform 1 0 33120 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1668240031
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1668240031
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_365
timestamp 1668240031
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_377
timestamp 1668240031
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_389
timestamp 1668240031
transform 1 0 36892 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_393
timestamp 1668240031
transform 1 0 37260 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1668240031
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1668240031
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1668240031
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1668240031
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1668240031
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1668240031
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_57
timestamp 1668240031
transform 1 0 6348 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_61
timestamp 1668240031
transform 1 0 6716 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_71
timestamp 1668240031
transform 1 0 7636 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_84
timestamp 1668240031
transform 1 0 8832 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_97
timestamp 1668240031
transform 1 0 10028 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_110
timestamp 1668240031
transform 1 0 11224 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_113
timestamp 1668240031
transform 1 0 11500 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_123
timestamp 1668240031
transform 1 0 12420 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_136
timestamp 1668240031
transform 1 0 13616 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_150
timestamp 1668240031
transform 1 0 14904 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_157
timestamp 1668240031
transform 1 0 15548 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_51_166
timestamp 1668240031
transform 1 0 16376 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_169
timestamp 1668240031
transform 1 0 16652 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_180
timestamp 1668240031
transform 1 0 17664 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_190
timestamp 1668240031
transform 1 0 18584 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_194
timestamp 1668240031
transform 1 0 18952 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_215
timestamp 1668240031
transform 1 0 20884 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_222
timestamp 1668240031
transform 1 0 21528 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_225
timestamp 1668240031
transform 1 0 21804 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_233
timestamp 1668240031
transform 1 0 22540 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_241
timestamp 1668240031
transform 1 0 23276 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_252
timestamp 1668240031
transform 1 0 24288 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_265
timestamp 1668240031
transform 1 0 25484 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_275
timestamp 1668240031
transform 1 0 26404 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1668240031
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_51_281
timestamp 1668240031
transform 1 0 26956 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_292
timestamp 1668240031
transform 1 0 27968 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_304
timestamp 1668240031
transform 1 0 29072 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_313
timestamp 1668240031
transform 1 0 29900 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_51_326
timestamp 1668240031
transform 1 0 31096 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_51_333
timestamp 1668240031
transform 1 0 31740 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_51_337
timestamp 1668240031
transform 1 0 32108 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_51_345
timestamp 1668240031
transform 1 0 32844 0 -1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_51_367
timestamp 1668240031
transform 1 0 34868 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_379
timestamp 1668240031
transform 1 0 35972 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1668240031
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_51_393
timestamp 1668240031
transform 1 0 37260 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1668240031
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1668240031
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1668240031
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1668240031
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1668240031
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_53
timestamp 1668240031
transform 1 0 5980 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_57
timestamp 1668240031
transform 1 0 6348 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_78
timestamp 1668240031
transform 1 0 8280 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_52_85
timestamp 1668240031
transform 1 0 8924 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_91
timestamp 1668240031
transform 1 0 9476 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_106
timestamp 1668240031
transform 1 0 10856 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_114
timestamp 1668240031
transform 1 0 11592 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_52_125
timestamp 1668240031
transform 1 0 12604 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_131
timestamp 1668240031
transform 1 0 13156 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_138
timestamp 1668240031
transform 1 0 13800 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_52_141
timestamp 1668240031
transform 1 0 14076 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_147
timestamp 1668240031
transform 1 0 14628 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_157
timestamp 1668240031
transform 1 0 15548 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_181
timestamp 1668240031
transform 1 0 17756 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_187
timestamp 1668240031
transform 1 0 18308 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_194
timestamp 1668240031
transform 1 0 18952 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_197
timestamp 1668240031
transform 1 0 19228 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_208
timestamp 1668240031
transform 1 0 20240 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_216
timestamp 1668240031
transform 1 0 20976 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_238
timestamp 1668240031
transform 1 0 23000 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_245
timestamp 1668240031
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1668240031
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_253
timestamp 1668240031
transform 1 0 24380 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_264
timestamp 1668240031
transform 1 0 25392 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_271
timestamp 1668240031
transform 1 0 26036 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_278
timestamp 1668240031
transform 1 0 26680 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_284
timestamp 1668240031
transform 1 0 27232 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_293
timestamp 1668240031
transform 1 0 28060 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_303
timestamp 1668240031
transform 1 0 28980 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1668240031
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_309
timestamp 1668240031
transform 1 0 29532 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_52_317
timestamp 1668240031
transform 1 0 30268 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_323
timestamp 1668240031
transform 1 0 30820 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_344
timestamp 1668240031
transform 1 0 32752 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_352
timestamp 1668240031
transform 1 0 33488 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_362
timestamp 1668240031
transform 1 0 34408 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_365
timestamp 1668240031
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_377
timestamp 1668240031
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_389
timestamp 1668240031
transform 1 0 36892 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_393
timestamp 1668240031
transform 1 0 37260 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1668240031
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1668240031
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1668240031
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_39
timestamp 1668240031
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1668240031
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1668240031
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_57
timestamp 1668240031
transform 1 0 6348 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_63
timestamp 1668240031
transform 1 0 6900 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_67
timestamp 1668240031
transform 1 0 7268 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_91
timestamp 1668240031
transform 1 0 9476 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_99
timestamp 1668240031
transform 1 0 10212 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_110
timestamp 1668240031
transform 1 0 11224 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_113
timestamp 1668240031
transform 1 0 11500 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_118
timestamp 1668240031
transform 1 0 11960 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_133
timestamp 1668240031
transform 1 0 13340 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_139
timestamp 1668240031
transform 1 0 13892 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_160
timestamp 1668240031
transform 1 0 15824 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_169
timestamp 1668240031
transform 1 0 16652 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_174
timestamp 1668240031
transform 1 0 17112 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_187
timestamp 1668240031
transform 1 0 18308 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_200
timestamp 1668240031
transform 1 0 19504 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_208
timestamp 1668240031
transform 1 0 20240 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_215
timestamp 1668240031
transform 1 0 20884 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_222
timestamp 1668240031
transform 1 0 21528 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_53_225
timestamp 1668240031
transform 1 0 21804 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_231
timestamp 1668240031
transform 1 0 22356 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_241
timestamp 1668240031
transform 1 0 23276 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_53_252
timestamp 1668240031
transform 1 0 24288 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_276
timestamp 1668240031
transform 1 0 26496 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_281
timestamp 1668240031
transform 1 0 26956 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_53_293
timestamp 1668240031
transform 1 0 28060 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_319
timestamp 1668240031
transform 1 0 30452 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_328
timestamp 1668240031
transform 1 0 31280 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_337
timestamp 1668240031
transform 1 0 32108 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_348
timestamp 1668240031
transform 1 0 33120 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_352
timestamp 1668240031
transform 1 0 33488 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_356
timestamp 1668240031
transform 1 0 33856 0 -1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_53_365
timestamp 1668240031
transform 1 0 34684 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_377
timestamp 1668240031
transform 1 0 35788 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_389
timestamp 1668240031
transform 1 0 36892 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_53_393
timestamp 1668240031
transform 1 0 37260 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_3
timestamp 1668240031
transform 1 0 1380 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_8
timestamp 1668240031
transform 1 0 1840 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_20
timestamp 1668240031
transform 1 0 2944 0 1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1668240031
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1668240031
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_53
timestamp 1668240031
transform 1 0 5980 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_62
timestamp 1668240031
transform 1 0 6808 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_69
timestamp 1668240031
transform 1 0 7452 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_82
timestamp 1668240031
transform 1 0 8648 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_85
timestamp 1668240031
transform 1 0 8924 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_90
timestamp 1668240031
transform 1 0 9384 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_114
timestamp 1668240031
transform 1 0 11592 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_138
timestamp 1668240031
transform 1 0 13800 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_141
timestamp 1668240031
transform 1 0 14076 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_152
timestamp 1668240031
transform 1 0 15088 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_156
timestamp 1668240031
transform 1 0 15456 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_166
timestamp 1668240031
transform 1 0 16376 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_194
timestamp 1668240031
transform 1 0 18952 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_197
timestamp 1668240031
transform 1 0 19228 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_202
timestamp 1668240031
transform 1 0 19688 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_209
timestamp 1668240031
transform 1 0 20332 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_233
timestamp 1668240031
transform 1 0 22540 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_246
timestamp 1668240031
transform 1 0 23736 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_54_253
timestamp 1668240031
transform 1 0 24380 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_276
timestamp 1668240031
transform 1 0 26496 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_283
timestamp 1668240031
transform 1 0 27140 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_287
timestamp 1668240031
transform 1 0 27508 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_294
timestamp 1668240031
transform 1 0 28152 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_306
timestamp 1668240031
transform 1 0 29256 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_309
timestamp 1668240031
transform 1 0 29532 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_317
timestamp 1668240031
transform 1 0 30268 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_324
timestamp 1668240031
transform 1 0 30912 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_349
timestamp 1668240031
transform 1 0 33212 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_356
timestamp 1668240031
transform 1 0 33856 0 1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_54_365
timestamp 1668240031
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_377
timestamp 1668240031
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_392
timestamp 1668240031
transform 1 0 37168 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1668240031
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1668240031
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_27
timestamp 1668240031
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_39
timestamp 1668240031
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1668240031
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1668240031
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_57
timestamp 1668240031
transform 1 0 6348 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_62
timestamp 1668240031
transform 1 0 6808 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_69
timestamp 1668240031
transform 1 0 7452 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_76
timestamp 1668240031
transform 1 0 8096 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_83
timestamp 1668240031
transform 1 0 8740 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_90
timestamp 1668240031
transform 1 0 9384 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_98
timestamp 1668240031
transform 1 0 10120 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_103
timestamp 1668240031
transform 1 0 10580 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_110
timestamp 1668240031
transform 1 0 11224 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_113
timestamp 1668240031
transform 1 0 11500 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_124
timestamp 1668240031
transform 1 0 12512 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_132
timestamp 1668240031
transform 1 0 13248 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_136
timestamp 1668240031
transform 1 0 13616 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_140
timestamp 1668240031
transform 1 0 13984 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1668240031
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1668240031
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_169
timestamp 1668240031
transform 1 0 16652 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_174
timestamp 1668240031
transform 1 0 17112 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_182
timestamp 1668240031
transform 1 0 17848 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_187
timestamp 1668240031
transform 1 0 18308 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_195
timestamp 1668240031
transform 1 0 19044 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_205
timestamp 1668240031
transform 1 0 19964 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_212
timestamp 1668240031
transform 1 0 20608 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_218
timestamp 1668240031
transform 1 0 21160 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_222
timestamp 1668240031
transform 1 0 21528 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_225
timestamp 1668240031
transform 1 0 21804 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_230
timestamp 1668240031
transform 1 0 22264 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_237
timestamp 1668240031
transform 1 0 22908 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_250
timestamp 1668240031
transform 1 0 24104 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_263
timestamp 1668240031
transform 1 0 25300 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_270
timestamp 1668240031
transform 1 0 25944 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_55_277
timestamp 1668240031
transform 1 0 26588 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_55_281
timestamp 1668240031
transform 1 0 26956 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_286
timestamp 1668240031
transform 1 0 27416 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_296
timestamp 1668240031
transform 1 0 28336 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_306
timestamp 1668240031
transform 1 0 29256 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_316
timestamp 1668240031
transform 1 0 30176 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_324
timestamp 1668240031
transform 1 0 30912 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_55_330
timestamp 1668240031
transform 1 0 31464 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_55_337
timestamp 1668240031
transform 1 0 32108 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_342
timestamp 1668240031
transform 1 0 32568 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_349
timestamp 1668240031
transform 1 0 33212 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_356
timestamp 1668240031
transform 1 0 33856 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_363
timestamp 1668240031
transform 1 0 34500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_375
timestamp 1668240031
transform 1 0 35604 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_387
timestamp 1668240031
transform 1 0 36708 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1668240031
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_55_393
timestamp 1668240031
transform 1 0 37260 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1668240031
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1668240031
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1668240031
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1668240031
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1668240031
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_53
timestamp 1668240031
transform 1 0 5980 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_81
timestamp 1668240031
transform 1 0 8556 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_56_85
timestamp 1668240031
transform 1 0 8924 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_91
timestamp 1668240031
transform 1 0 9476 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_101
timestamp 1668240031
transform 1 0 10396 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_110
timestamp 1668240031
transform 1 0 11224 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_123
timestamp 1668240031
transform 1 0 12420 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_129
timestamp 1668240031
transform 1 0 12972 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1668240031
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1668240031
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_141
timestamp 1668240031
transform 1 0 14076 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_156
timestamp 1668240031
transform 1 0 15456 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_181
timestamp 1668240031
transform 1 0 17756 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_194
timestamp 1668240031
transform 1 0 18952 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_197
timestamp 1668240031
transform 1 0 19228 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_56_219
timestamp 1668240031
transform 1 0 21252 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_236
timestamp 1668240031
transform 1 0 22816 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_56_249
timestamp 1668240031
transform 1 0 24012 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_56_253
timestamp 1668240031
transform 1 0 24380 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_56_264
timestamp 1668240031
transform 1 0 25392 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_273
timestamp 1668240031
transform 1 0 26220 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_280
timestamp 1668240031
transform 1 0 26864 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_292
timestamp 1668240031
transform 1 0 27968 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_303
timestamp 1668240031
transform 1 0 28980 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1668240031
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_309
timestamp 1668240031
transform 1 0 29532 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_320
timestamp 1668240031
transform 1 0 30544 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_324
timestamp 1668240031
transform 1 0 30912 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_345
timestamp 1668240031
transform 1 0 32844 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_362
timestamp 1668240031
transform 1 0 34408 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 1668240031
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_377
timestamp 1668240031
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_389
timestamp 1668240031
transform 1 0 36892 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_393
timestamp 1668240031
transform 1 0 37260 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1668240031
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1668240031
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1668240031
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 1668240031
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1668240031
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1668240031
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_57
timestamp 1668240031
transform 1 0 6348 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_65
timestamp 1668240031
transform 1 0 7084 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_69
timestamp 1668240031
transform 1 0 7452 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_93
timestamp 1668240031
transform 1 0 9660 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_106
timestamp 1668240031
transform 1 0 10856 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_57_113
timestamp 1668240031
transform 1 0 11500 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_57_141
timestamp 1668240031
transform 1 0 14076 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_149
timestamp 1668240031
transform 1 0 14812 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_153
timestamp 1668240031
transform 1 0 15180 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_166
timestamp 1668240031
transform 1 0 16376 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_57_169
timestamp 1668240031
transform 1 0 16652 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_175
timestamp 1668240031
transform 1 0 17204 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_196
timestamp 1668240031
transform 1 0 19136 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_211
timestamp 1668240031
transform 1 0 20516 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1668240031
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_225
timestamp 1668240031
transform 1 0 21804 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_247
timestamp 1668240031
transform 1 0 23828 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_254
timestamp 1668240031
transform 1 0 24472 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_278
timestamp 1668240031
transform 1 0 26680 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1668240031
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_299
timestamp 1668240031
transform 1 0 28612 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_308
timestamp 1668240031
transform 1 0 29440 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_323
timestamp 1668240031
transform 1 0 30820 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_330
timestamp 1668240031
transform 1 0 31464 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_57_337
timestamp 1668240031
transform 1 0 32108 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_342
timestamp 1668240031
transform 1 0 32568 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_349
timestamp 1668240031
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_361
timestamp 1668240031
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_373
timestamp 1668240031
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1668240031
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1668240031
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_57_393
timestamp 1668240031
transform 1 0 37260 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1668240031
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1668240031
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1668240031
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1668240031
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1668240031
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1668240031
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_65
timestamp 1668240031
transform 1 0 7084 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_82
timestamp 1668240031
transform 1 0 8648 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_85
timestamp 1668240031
transform 1 0 8924 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_96
timestamp 1668240031
transform 1 0 9936 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_100
timestamp 1668240031
transform 1 0 10304 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_121
timestamp 1668240031
transform 1 0 12236 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_134
timestamp 1668240031
transform 1 0 13432 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_58_141
timestamp 1668240031
transform 1 0 14076 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_152
timestamp 1668240031
transform 1 0 15088 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_156
timestamp 1668240031
transform 1 0 15456 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_166
timestamp 1668240031
transform 1 0 16376 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_173
timestamp 1668240031
transform 1 0 17020 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_180
timestamp 1668240031
transform 1 0 17664 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_187
timestamp 1668240031
transform 1 0 18308 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_194
timestamp 1668240031
transform 1 0 18952 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_58_197
timestamp 1668240031
transform 1 0 19228 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_209
timestamp 1668240031
transform 1 0 20332 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_216
timestamp 1668240031
transform 1 0 20976 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_228
timestamp 1668240031
transform 1 0 22080 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_232
timestamp 1668240031
transform 1 0 22448 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1668240031
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1668240031
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_253
timestamp 1668240031
transform 1 0 24380 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_58_279
timestamp 1668240031
transform 1 0 26772 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_287
timestamp 1668240031
transform 1 0 27508 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_58_297
timestamp 1668240031
transform 1 0 28428 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_305
timestamp 1668240031
transform 1 0 29164 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_58_309
timestamp 1668240031
transform 1 0 29532 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_58_314
timestamp 1668240031
transform 1 0 29992 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_322
timestamp 1668240031
transform 1 0 30728 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_343
timestamp 1668240031
transform 1 0 32660 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_350
timestamp 1668240031
transform 1 0 33304 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_362
timestamp 1668240031
transform 1 0 34408 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_365
timestamp 1668240031
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_377
timestamp 1668240031
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_389
timestamp 1668240031
transform 1 0 36892 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_393
timestamp 1668240031
transform 1 0 37260 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1668240031
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1668240031
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 1668240031
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_39
timestamp 1668240031
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1668240031
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1668240031
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1668240031
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_69
timestamp 1668240031
transform 1 0 7452 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_77
timestamp 1668240031
transform 1 0 8188 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_59_89
timestamp 1668240031
transform 1 0 9292 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_97
timestamp 1668240031
transform 1 0 10028 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_59_103
timestamp 1668240031
transform 1 0 10580 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_110
timestamp 1668240031
transform 1 0 11224 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_113
timestamp 1668240031
transform 1 0 11500 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_124
timestamp 1668240031
transform 1 0 12512 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_128
timestamp 1668240031
transform 1 0 12880 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_149
timestamp 1668240031
transform 1 0 14812 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_155
timestamp 1668240031
transform 1 0 15364 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_159
timestamp 1668240031
transform 1 0 15732 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_166
timestamp 1668240031
transform 1 0 16376 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_59_169
timestamp 1668240031
transform 1 0 16652 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_59_180
timestamp 1668240031
transform 1 0 17664 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_193
timestamp 1668240031
transform 1 0 18860 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_59_219
timestamp 1668240031
transform 1 0 21252 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1668240031
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_225
timestamp 1668240031
transform 1 0 21804 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_249
timestamp 1668240031
transform 1 0 24012 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_262
timestamp 1668240031
transform 1 0 25208 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_269
timestamp 1668240031
transform 1 0 25852 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_276
timestamp 1668240031
transform 1 0 26496 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_281
timestamp 1668240031
transform 1 0 26956 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_289
timestamp 1668240031
transform 1 0 27692 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_300
timestamp 1668240031
transform 1 0 28704 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_307
timestamp 1668240031
transform 1 0 29348 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_318
timestamp 1668240031
transform 1 0 30360 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_326
timestamp 1668240031
transform 1 0 31096 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_59_333
timestamp 1668240031
transform 1 0 31740 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_59_337
timestamp 1668240031
transform 1 0 32108 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_359
timestamp 1668240031
transform 1 0 34132 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_371
timestamp 1668240031
transform 1 0 35236 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_383
timestamp 1668240031
transform 1 0 36340 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1668240031
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_59_393
timestamp 1668240031
transform 1 0 37260 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_3
timestamp 1668240031
transform 1 0 1380 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_8
timestamp 1668240031
transform 1 0 1840 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_20
timestamp 1668240031
transform 1 0 2944 0 1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1668240031
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1668240031
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_53
timestamp 1668240031
transform 1 0 5980 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_59
timestamp 1668240031
transform 1 0 6532 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_80
timestamp 1668240031
transform 1 0 8464 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_85
timestamp 1668240031
transform 1 0 8924 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_96
timestamp 1668240031
transform 1 0 9936 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_109
timestamp 1668240031
transform 1 0 11132 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_113
timestamp 1668240031
transform 1 0 11500 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_117
timestamp 1668240031
transform 1 0 11868 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_124
timestamp 1668240031
transform 1 0 12512 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_131
timestamp 1668240031
transform 1 0 13156 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_138
timestamp 1668240031
transform 1 0 13800 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_141
timestamp 1668240031
transform 1 0 14076 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_163
timestamp 1668240031
transform 1 0 16100 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_187
timestamp 1668240031
transform 1 0 18308 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_194
timestamp 1668240031
transform 1 0 18952 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_197
timestamp 1668240031
transform 1 0 19228 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_208
timestamp 1668240031
transform 1 0 20240 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_232
timestamp 1668240031
transform 1 0 22448 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_240
timestamp 1668240031
transform 1 0 23184 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_250
timestamp 1668240031
transform 1 0 24104 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_253
timestamp 1668240031
transform 1 0 24380 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_264
timestamp 1668240031
transform 1 0 25392 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_277
timestamp 1668240031
transform 1 0 26588 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_287
timestamp 1668240031
transform 1 0 27508 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_300
timestamp 1668240031
transform 1 0 28704 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_309
timestamp 1668240031
transform 1 0 29532 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_60_317
timestamp 1668240031
transform 1 0 30268 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_325
timestamp 1668240031
transform 1 0 31004 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_347
timestamp 1668240031
transform 1 0 33028 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_354
timestamp 1668240031
transform 1 0 33672 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_362
timestamp 1668240031
transform 1 0 34408 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1668240031
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_377
timestamp 1668240031
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_392
timestamp 1668240031
transform 1 0 37168 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1668240031
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1668240031
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1668240031
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_39
timestamp 1668240031
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1668240031
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1668240031
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_57
timestamp 1668240031
transform 1 0 6348 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_62
timestamp 1668240031
transform 1 0 6808 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_69
timestamp 1668240031
transform 1 0 7452 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_93
timestamp 1668240031
transform 1 0 9660 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_110
timestamp 1668240031
transform 1 0 11224 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_113
timestamp 1668240031
transform 1 0 11500 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_124
timestamp 1668240031
transform 1 0 12512 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_137
timestamp 1668240031
transform 1 0 13708 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_61_146
timestamp 1668240031
transform 1 0 14536 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_159
timestamp 1668240031
transform 1 0 15732 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_166
timestamp 1668240031
transform 1 0 16376 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_169
timestamp 1668240031
transform 1 0 16652 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_177
timestamp 1668240031
transform 1 0 17388 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_187
timestamp 1668240031
transform 1 0 18308 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_61_198
timestamp 1668240031
transform 1 0 19320 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_202
timestamp 1668240031
transform 1 0 19688 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_212
timestamp 1668240031
transform 1 0 20608 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_219
timestamp 1668240031
transform 1 0 21252 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1668240031
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_225
timestamp 1668240031
transform 1 0 21804 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_230
timestamp 1668240031
transform 1 0 22264 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_234
timestamp 1668240031
transform 1 0 22632 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_238
timestamp 1668240031
transform 1 0 23000 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_242
timestamp 1668240031
transform 1 0 23368 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_252
timestamp 1668240031
transform 1 0 24288 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_61_278
timestamp 1668240031
transform 1 0 26680 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_281
timestamp 1668240031
transform 1 0 26956 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_61_297
timestamp 1668240031
transform 1 0 28428 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_307
timestamp 1668240031
transform 1 0 29348 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_311
timestamp 1668240031
transform 1 0 29716 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_317
timestamp 1668240031
transform 1 0 30268 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_326
timestamp 1668240031
transform 1 0 31096 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_61_333
timestamp 1668240031
transform 1 0 31740 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_61_337
timestamp 1668240031
transform 1 0 32108 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_359
timestamp 1668240031
transform 1 0 34132 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_371
timestamp 1668240031
transform 1 0 35236 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_383
timestamp 1668240031
transform 1 0 36340 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1668240031
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_61_393
timestamp 1668240031
transform 1 0 37260 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1668240031
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1668240031
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1668240031
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1668240031
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1668240031
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1668240031
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_65
timestamp 1668240031
transform 1 0 7084 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_69
timestamp 1668240031
transform 1 0 7452 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_82
timestamp 1668240031
transform 1 0 8648 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_62_85
timestamp 1668240031
transform 1 0 8924 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_91
timestamp 1668240031
transform 1 0 9476 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_101
timestamp 1668240031
transform 1 0 10396 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_125
timestamp 1668240031
transform 1 0 12604 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_138
timestamp 1668240031
transform 1 0 13800 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_62_141
timestamp 1668240031
transform 1 0 14076 0 1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_62_158
timestamp 1668240031
transform 1 0 15640 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_170
timestamp 1668240031
transform 1 0 16744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_174
timestamp 1668240031
transform 1 0 17112 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_181
timestamp 1668240031
transform 1 0 17756 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_194
timestamp 1668240031
transform 1 0 18952 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_197
timestamp 1668240031
transform 1 0 19228 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_201
timestamp 1668240031
transform 1 0 19596 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_211
timestamp 1668240031
transform 1 0 20516 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_223
timestamp 1668240031
transform 1 0 21620 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_62_228
timestamp 1668240031
transform 1 0 22080 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_236
timestamp 1668240031
transform 1 0 22816 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_247
timestamp 1668240031
transform 1 0 23828 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1668240031
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_253
timestamp 1668240031
transform 1 0 24380 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_264
timestamp 1668240031
transform 1 0 25392 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_271
timestamp 1668240031
transform 1 0 26036 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_278
timestamp 1668240031
transform 1 0 26680 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_286
timestamp 1668240031
transform 1 0 27416 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_294
timestamp 1668240031
transform 1 0 28152 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_304
timestamp 1668240031
transform 1 0 29072 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_309
timestamp 1668240031
transform 1 0 29532 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_317
timestamp 1668240031
transform 1 0 30268 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_324
timestamp 1668240031
transform 1 0 30912 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_348
timestamp 1668240031
transform 1 0 33120 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_355
timestamp 1668240031
transform 1 0 33764 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1668240031
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_365
timestamp 1668240031
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_377
timestamp 1668240031
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_389
timestamp 1668240031
transform 1 0 36892 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_393
timestamp 1668240031
transform 1 0 37260 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1668240031
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 1668240031
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_27
timestamp 1668240031
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_39
timestamp 1668240031
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1668240031
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1668240031
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1668240031
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 1668240031
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_81
timestamp 1668240031
transform 1 0 8556 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_85
timestamp 1668240031
transform 1 0 8924 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_89
timestamp 1668240031
transform 1 0 9292 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_93
timestamp 1668240031
transform 1 0 9660 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_103
timestamp 1668240031
transform 1 0 10580 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_110
timestamp 1668240031
transform 1 0 11224 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_113
timestamp 1668240031
transform 1 0 11500 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_120
timestamp 1668240031
transform 1 0 12144 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_124
timestamp 1668240031
transform 1 0 12512 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_134
timestamp 1668240031
transform 1 0 13432 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_158
timestamp 1668240031
transform 1 0 15640 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_162
timestamp 1668240031
transform 1 0 16008 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_166
timestamp 1668240031
transform 1 0 16376 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_63_169
timestamp 1668240031
transform 1 0 16652 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_181
timestamp 1668240031
transform 1 0 17756 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_205
timestamp 1668240031
transform 1 0 19964 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_212
timestamp 1668240031
transform 1 0 20608 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_218
timestamp 1668240031
transform 1 0 21160 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_222
timestamp 1668240031
transform 1 0 21528 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_63_225
timestamp 1668240031
transform 1 0 21804 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_248
timestamp 1668240031
transform 1 0 23920 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_261
timestamp 1668240031
transform 1 0 25116 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_274
timestamp 1668240031
transform 1 0 26312 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_63_281
timestamp 1668240031
transform 1 0 26956 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_63_286
timestamp 1668240031
transform 1 0 27416 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_298
timestamp 1668240031
transform 1 0 28520 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_306
timestamp 1668240031
transform 1 0 29256 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_317
timestamp 1668240031
transform 1 0 30268 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_324
timestamp 1668240031
transform 1 0 30912 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_337
timestamp 1668240031
transform 1 0 32108 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_359
timestamp 1668240031
transform 1 0 34132 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_371
timestamp 1668240031
transform 1 0 35236 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_383
timestamp 1668240031
transform 1 0 36340 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1668240031
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_63_393
timestamp 1668240031
transform 1 0 37260 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_3
timestamp 1668240031
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_15
timestamp 1668240031
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1668240031
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1668240031
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_41
timestamp 1668240031
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_53
timestamp 1668240031
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_65
timestamp 1668240031
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_77
timestamp 1668240031
transform 1 0 8188 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_82
timestamp 1668240031
transform 1 0 8648 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_85
timestamp 1668240031
transform 1 0 8924 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_107
timestamp 1668240031
transform 1 0 10948 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_64_135
timestamp 1668240031
transform 1 0 13524 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1668240031
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_141
timestamp 1668240031
transform 1 0 14076 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_145
timestamp 1668240031
transform 1 0 14444 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_155
timestamp 1668240031
transform 1 0 15364 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_179
timestamp 1668240031
transform 1 0 17572 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_64_194
timestamp 1668240031
transform 1 0 18952 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_197
timestamp 1668240031
transform 1 0 19228 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_204
timestamp 1668240031
transform 1 0 19872 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_228
timestamp 1668240031
transform 1 0 22080 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_232
timestamp 1668240031
transform 1 0 22448 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_236
timestamp 1668240031
transform 1 0 22816 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_240
timestamp 1668240031
transform 1 0 23184 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_250
timestamp 1668240031
transform 1 0 24104 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_253
timestamp 1668240031
transform 1 0 24380 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_64_279
timestamp 1668240031
transform 1 0 26772 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_287
timestamp 1668240031
transform 1 0 27508 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_296
timestamp 1668240031
transform 1 0 28336 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_306
timestamp 1668240031
transform 1 0 29256 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_309
timestamp 1668240031
transform 1 0 29532 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_318
timestamp 1668240031
transform 1 0 30360 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_324
timestamp 1668240031
transform 1 0 30912 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_346
timestamp 1668240031
transform 1 0 32936 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_353
timestamp 1668240031
transform 1 0 33580 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_361
timestamp 1668240031
transform 1 0 34316 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_365
timestamp 1668240031
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_377
timestamp 1668240031
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_389
timestamp 1668240031
transform 1 0 36892 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_393
timestamp 1668240031
transform 1 0 37260 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_3
timestamp 1668240031
transform 1 0 1380 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_65_8
timestamp 1668240031
transform 1 0 1840 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_20
timestamp 1668240031
transform 1 0 2944 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_32
timestamp 1668240031
transform 1 0 4048 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_65_40
timestamp 1668240031
transform 1 0 4784 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_65_46
timestamp 1668240031
transform 1 0 5336 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_65_54
timestamp 1668240031
transform 1 0 6072 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_65_57
timestamp 1668240031
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_69
timestamp 1668240031
transform 1 0 7452 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_75
timestamp 1668240031
transform 1 0 8004 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_79
timestamp 1668240031
transform 1 0 8372 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_65_87
timestamp 1668240031
transform 1 0 9108 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_65_93
timestamp 1668240031
transform 1 0 9660 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_97
timestamp 1668240031
transform 1 0 10028 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_101
timestamp 1668240031
transform 1 0 10396 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_108
timestamp 1668240031
transform 1 0 11040 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_65_113
timestamp 1668240031
transform 1 0 11500 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_65_119
timestamp 1668240031
transform 1 0 12052 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_65_132
timestamp 1668240031
transform 1 0 13248 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_138
timestamp 1668240031
transform 1 0 13800 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_148
timestamp 1668240031
transform 1 0 14720 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_156
timestamp 1668240031
transform 1 0 15456 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_160
timestamp 1668240031
transform 1 0 15824 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_65_169
timestamp 1668240031
transform 1 0 16652 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_191
timestamp 1668240031
transform 1 0 18676 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_198
timestamp 1668240031
transform 1 0 19320 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_211
timestamp 1668240031
transform 1 0 20516 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_65_218
timestamp 1668240031
transform 1 0 21160 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_65_225
timestamp 1668240031
transform 1 0 21804 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_247
timestamp 1668240031
transform 1 0 23828 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_271
timestamp 1668240031
transform 1 0 26036 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_278
timestamp 1668240031
transform 1 0 26680 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_65_281
timestamp 1668240031
transform 1 0 26956 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_65_290
timestamp 1668240031
transform 1 0 27784 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_300
timestamp 1668240031
transform 1 0 28704 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_310
timestamp 1668240031
transform 1 0 29624 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_334
timestamp 1668240031
transform 1 0 31832 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_337
timestamp 1668240031
transform 1 0 32108 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_359
timestamp 1668240031
transform 1 0 34132 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_65_366
timestamp 1668240031
transform 1 0 34776 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_378
timestamp 1668240031
transform 1 0 35880 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_65_390
timestamp 1668240031
transform 1 0 36984 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_65_393
timestamp 1668240031
transform 1 0 37260 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_3
timestamp 1668240031
transform 1 0 1380 0 1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_66_10
timestamp 1668240031
transform 1 0 2024 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_22
timestamp 1668240031
transform 1 0 3128 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_66_29
timestamp 1668240031
transform 1 0 3772 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_37
timestamp 1668240031
transform 1 0 4508 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_66_42
timestamp 1668240031
transform 1 0 4968 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_66_54
timestamp 1668240031
transform 1 0 6072 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_66_57
timestamp 1668240031
transform 1 0 6348 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_66_69
timestamp 1668240031
transform 1 0 7452 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_66_74
timestamp 1668240031
transform 1 0 7912 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_82
timestamp 1668240031
transform 1 0 8648 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_66_85
timestamp 1668240031
transform 1 0 8924 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_66_96
timestamp 1668240031
transform 1 0 9936 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_103
timestamp 1668240031
transform 1 0 10580 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_110
timestamp 1668240031
transform 1 0 11224 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_66_113
timestamp 1668240031
transform 1 0 11500 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_66_124
timestamp 1668240031
transform 1 0 12512 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_131
timestamp 1668240031
transform 1 0 13156 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_138
timestamp 1668240031
transform 1 0 13800 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_141
timestamp 1668240031
transform 1 0 14076 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_148
timestamp 1668240031
transform 1 0 14720 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_66_155
timestamp 1668240031
transform 1 0 15364 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_166
timestamp 1668240031
transform 1 0 16376 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_169
timestamp 1668240031
transform 1 0 16652 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_173
timestamp 1668240031
transform 1 0 17020 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_177
timestamp 1668240031
transform 1 0 17388 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_66_190
timestamp 1668240031
transform 1 0 18584 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_66_197
timestamp 1668240031
transform 1 0 19228 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_208
timestamp 1668240031
transform 1 0 20240 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_66_221
timestamp 1668240031
transform 1 0 21436 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_66_225
timestamp 1668240031
transform 1 0 21804 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_66_234
timestamp 1668240031
transform 1 0 22632 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_241
timestamp 1668240031
transform 1 0 23276 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_248
timestamp 1668240031
transform 1 0 23920 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_253
timestamp 1668240031
transform 1 0 24380 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_258
timestamp 1668240031
transform 1 0 24840 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_265
timestamp 1668240031
transform 1 0 25484 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_66_272
timestamp 1668240031
transform 1 0 26128 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_66_281
timestamp 1668240031
transform 1 0 26956 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_66_293
timestamp 1668240031
transform 1 0 28060 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_66_302
timestamp 1668240031
transform 1 0 28888 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_66_309
timestamp 1668240031
transform 1 0 29532 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_316
timestamp 1668240031
transform 1 0 30176 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_323
timestamp 1668240031
transform 1 0 30820 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_66_330
timestamp 1668240031
transform 1 0 31464 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_66_337
timestamp 1668240031
transform 1 0 32108 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_342
timestamp 1668240031
transform 1 0 32568 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_66_349
timestamp 1668240031
transform 1 0 33212 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_357
timestamp 1668240031
transform 1 0 33948 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_362
timestamp 1668240031
transform 1 0 34408 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_66_365
timestamp 1668240031
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_377
timestamp 1668240031
transform 1 0 35788 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_385
timestamp 1668240031
transform 1 0 36524 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_390
timestamp 1668240031
transform 1 0 36984 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_66_393
timestamp 1668240031
transform 1 0 37260 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1668240031
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1668240031
transform -1 0 37628 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1668240031
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1668240031
transform -1 0 37628 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1668240031
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1668240031
transform -1 0 37628 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1668240031
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1668240031
transform -1 0 37628 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1668240031
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1668240031
transform -1 0 37628 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1668240031
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1668240031
transform -1 0 37628 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1668240031
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1668240031
transform -1 0 37628 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1668240031
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1668240031
transform -1 0 37628 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1668240031
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1668240031
transform -1 0 37628 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1668240031
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1668240031
transform -1 0 37628 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1668240031
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1668240031
transform -1 0 37628 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1668240031
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1668240031
transform -1 0 37628 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1668240031
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1668240031
transform -1 0 37628 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1668240031
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1668240031
transform -1 0 37628 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1668240031
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1668240031
transform -1 0 37628 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1668240031
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1668240031
transform -1 0 37628 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1668240031
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1668240031
transform -1 0 37628 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1668240031
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1668240031
transform -1 0 37628 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1668240031
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1668240031
transform -1 0 37628 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1668240031
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1668240031
transform -1 0 37628 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1668240031
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1668240031
transform -1 0 37628 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1668240031
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1668240031
transform -1 0 37628 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1668240031
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1668240031
transform -1 0 37628 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1668240031
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1668240031
transform -1 0 37628 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1668240031
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1668240031
transform -1 0 37628 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1668240031
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1668240031
transform -1 0 37628 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1668240031
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1668240031
transform -1 0 37628 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1668240031
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1668240031
transform -1 0 37628 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1668240031
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1668240031
transform -1 0 37628 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1668240031
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1668240031
transform -1 0 37628 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1668240031
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1668240031
transform -1 0 37628 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1668240031
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1668240031
transform -1 0 37628 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1668240031
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1668240031
transform -1 0 37628 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1668240031
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1668240031
transform -1 0 37628 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1668240031
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1668240031
transform -1 0 37628 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1668240031
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1668240031
transform -1 0 37628 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1668240031
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1668240031
transform -1 0 37628 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1668240031
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1668240031
transform -1 0 37628 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1668240031
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1668240031
transform -1 0 37628 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1668240031
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1668240031
transform -1 0 37628 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1668240031
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1668240031
transform -1 0 37628 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1668240031
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1668240031
transform -1 0 37628 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1668240031
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1668240031
transform -1 0 37628 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1668240031
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1668240031
transform -1 0 37628 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1668240031
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1668240031
transform -1 0 37628 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1668240031
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1668240031
transform -1 0 37628 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1668240031
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1668240031
transform -1 0 37628 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1668240031
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1668240031
transform -1 0 37628 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1668240031
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1668240031
transform -1 0 37628 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1668240031
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1668240031
transform -1 0 37628 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1668240031
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1668240031
transform -1 0 37628 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1668240031
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1668240031
transform -1 0 37628 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1668240031
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1668240031
transform -1 0 37628 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1668240031
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1668240031
transform -1 0 37628 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1668240031
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1668240031
transform -1 0 37628 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1668240031
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1668240031
transform -1 0 37628 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1668240031
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1668240031
transform -1 0 37628 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1668240031
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1668240031
transform -1 0 37628 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1668240031
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1668240031
transform -1 0 37628 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1668240031
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1668240031
transform -1 0 37628 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1668240031
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1668240031
transform -1 0 37628 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1668240031
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1668240031
transform -1 0 37628 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1668240031
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1668240031
transform -1 0 37628 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1668240031
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1668240031
transform -1 0 37628 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1668240031
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1668240031
transform -1 0 37628 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1668240031
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1668240031
transform -1 0 37628 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1668240031
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1668240031
transform -1 0 37628 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1668240031
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1668240031
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1668240031
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1668240031
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1668240031
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1668240031
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1668240031
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1668240031
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1668240031
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1668240031
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1668240031
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1668240031
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1668240031
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1668240031
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1668240031
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1668240031
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1668240031
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1668240031
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1668240031
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1668240031
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1668240031
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1668240031
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1668240031
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1668240031
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1668240031
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1668240031
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1668240031
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1668240031
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1668240031
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1668240031
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1668240031
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1668240031
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1668240031
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1668240031
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1668240031
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1668240031
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1668240031
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1668240031
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1668240031
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1668240031
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1668240031
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1668240031
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1668240031
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1668240031
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1668240031
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1668240031
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1668240031
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1668240031
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1668240031
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1668240031
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1668240031
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1668240031
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1668240031
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1668240031
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1668240031
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1668240031
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1668240031
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1668240031
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1668240031
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1668240031
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1668240031
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1668240031
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1668240031
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1668240031
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1668240031
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1668240031
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1668240031
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1668240031
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1668240031
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1668240031
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1668240031
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1668240031
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1668240031
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1668240031
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1668240031
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1668240031
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1668240031
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1668240031
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1668240031
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1668240031
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1668240031
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1668240031
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1668240031
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1668240031
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1668240031
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1668240031
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1668240031
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1668240031
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1668240031
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1668240031
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1668240031
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1668240031
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1668240031
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1668240031
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1668240031
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1668240031
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1668240031
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1668240031
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1668240031
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1668240031
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1668240031
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1668240031
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1668240031
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1668240031
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1668240031
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1668240031
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1668240031
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1668240031
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1668240031
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1668240031
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1668240031
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1668240031
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1668240031
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1668240031
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1668240031
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1668240031
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1668240031
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1668240031
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1668240031
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1668240031
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1668240031
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1668240031
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1668240031
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1668240031
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1668240031
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1668240031
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1668240031
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1668240031
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1668240031
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1668240031
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1668240031
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1668240031
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1668240031
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1668240031
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1668240031
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1668240031
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1668240031
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1668240031
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1668240031
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1668240031
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1668240031
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1668240031
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1668240031
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1668240031
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1668240031
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1668240031
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1668240031
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1668240031
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1668240031
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1668240031
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1668240031
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1668240031
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1668240031
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1668240031
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1668240031
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1668240031
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1668240031
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1668240031
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1668240031
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1668240031
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1668240031
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1668240031
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1668240031
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1668240031
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1668240031
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1668240031
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1668240031
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1668240031
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1668240031
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1668240031
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1668240031
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1668240031
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1668240031
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1668240031
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1668240031
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1668240031
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1668240031
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1668240031
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1668240031
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1668240031
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1668240031
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1668240031
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1668240031
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1668240031
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1668240031
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1668240031
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1668240031
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1668240031
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1668240031
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1668240031
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1668240031
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1668240031
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1668240031
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1668240031
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1668240031
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1668240031
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1668240031
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1668240031
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1668240031
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1668240031
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1668240031
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1668240031
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1668240031
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1668240031
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1668240031
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1668240031
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1668240031
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1668240031
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1668240031
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1668240031
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1668240031
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1668240031
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1668240031
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1668240031
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1668240031
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1668240031
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1668240031
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1668240031
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1668240031
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1668240031
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1668240031
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1668240031
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1668240031
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1668240031
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1668240031
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1668240031
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1668240031
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1668240031
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1668240031
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1668240031
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1668240031
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1668240031
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1668240031
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1668240031
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1668240031
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1668240031
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1668240031
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1668240031
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1668240031
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1668240031
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1668240031
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1668240031
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1668240031
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1668240031
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1668240031
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1668240031
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1668240031
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1668240031
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1668240031
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1668240031
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1668240031
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1668240031
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1668240031
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1668240031
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1668240031
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1668240031
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1668240031
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1668240031
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1668240031
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1668240031
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1668240031
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1668240031
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1668240031
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1668240031
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1668240031
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1668240031
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1668240031
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1668240031
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1668240031
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1668240031
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1668240031
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1668240031
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1668240031
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1668240031
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1668240031
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1668240031
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1668240031
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1668240031
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1668240031
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1668240031
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1668240031
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1668240031
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1668240031
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1668240031
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1668240031
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1668240031
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1668240031
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1668240031
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1668240031
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1668240031
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1668240031
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1668240031
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1668240031
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1668240031
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1668240031
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1668240031
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1668240031
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1668240031
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1668240031
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1668240031
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1668240031
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1668240031
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1668240031
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1668240031
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1668240031
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1668240031
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1668240031
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1668240031
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1668240031
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1668240031
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1668240031
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1668240031
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1668240031
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1668240031
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1668240031
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1668240031
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1668240031
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1668240031
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1668240031
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1668240031
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1668240031
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1668240031
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1668240031
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1668240031
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1668240031
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1668240031
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1668240031
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1668240031
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1668240031
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1668240031
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1668240031
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1668240031
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1668240031
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1668240031
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1668240031
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1668240031
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1668240031
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1668240031
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1668240031
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1668240031
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1668240031
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1668240031
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1668240031
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1668240031
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1668240031
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1668240031
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1668240031
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1668240031
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1668240031
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1668240031
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1668240031
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1668240031
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1668240031
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1668240031
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1668240031
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1668240031
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1668240031
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1668240031
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1668240031
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1668240031
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1668240031
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1668240031
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1668240031
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1668240031
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1668240031
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1668240031
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1668240031
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1668240031
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1668240031
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1668240031
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1668240031
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1668240031
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1668240031
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1668240031
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1668240031
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1668240031
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1668240031
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1668240031
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1668240031
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1668240031
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1668240031
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1668240031
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1668240031
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1668240031
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1668240031
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1668240031
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1668240031
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1668240031
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1668240031
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1668240031
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1668240031
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1668240031
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1668240031
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1668240031
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1668240031
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1668240031
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1668240031
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1668240031
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1668240031
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1668240031
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1668240031
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1668240031
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1668240031
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1668240031
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1668240031
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1668240031
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1668240031
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1668240031
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1668240031
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1668240031
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1668240031
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1668240031
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1668240031
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1668240031
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1668240031
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1668240031
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1668240031
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1668240031
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1668240031
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1668240031
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1668240031
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1668240031
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1668240031
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1668240031
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1668240031
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1668240031
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1668240031
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1668240031
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1668240031
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1668240031
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1668240031
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1668240031
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1668240031
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1668240031
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1668240031
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1668240031
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1668240031
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1668240031
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1668240031
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1668240031
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1668240031
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1668240031
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1668240031
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1668240031
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1668240031
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1668240031
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1668240031
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1668240031
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1668240031
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1668240031
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1668240031
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1668240031
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1668240031
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1668240031
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1668240031
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1668240031
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1668240031
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1668240031
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1668240031
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1668240031
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1668240031
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1668240031
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1668240031
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1668240031
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1668240031
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1668240031
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1668240031
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1668240031
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1668240031
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1668240031
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1668240031
transform 1 0 6256 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1668240031
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1668240031
transform 1 0 11408 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1668240031
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1668240031
transform 1 0 16560 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1668240031
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1668240031
transform 1 0 21712 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1668240031
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1668240031
transform 1 0 26864 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1668240031
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1668240031
transform 1 0 32016 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1668240031
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1668240031
transform 1 0 37168 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  _0992_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1668240031
transform 1 0 27140 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0993_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1668240031
transform 1 0 30912 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0994_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1668240031
transform -1 0 31740 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0995_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1668240031
transform 1 0 31556 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0996_
timestamp 1668240031
transform 1 0 27232 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0997_
timestamp 1668240031
transform 1 0 26404 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0998_
timestamp 1668240031
transform 1 0 28336 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0999_
timestamp 1668240031
transform 1 0 27140 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1000_
timestamp 1668240031
transform -1 0 30636 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1001_
timestamp 1668240031
transform 1 0 30820 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1002_
timestamp 1668240031
transform -1 0 33304 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1003_
timestamp 1668240031
transform -1 0 33120 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1004_
timestamp 1668240031
transform 1 0 32936 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1005_
timestamp 1668240031
transform -1 0 32568 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1006_
timestamp 1668240031
transform -1 0 33396 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1007_
timestamp 1668240031
transform 1 0 33948 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1008_
timestamp 1668240031
transform -1 0 34040 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1009_
timestamp 1668240031
transform 1 0 33948 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1010_
timestamp 1668240031
transform -1 0 33948 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1011_
timestamp 1668240031
transform 1 0 34868 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1012_
timestamp 1668240031
transform 1 0 29440 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1013_
timestamp 1668240031
transform -1 0 28796 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1014_
timestamp 1668240031
transform 1 0 22632 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1015_
timestamp 1668240031
transform -1 0 23644 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1016_
timestamp 1668240031
transform -1 0 24840 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1017_
timestamp 1668240031
transform 1 0 20056 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1018_
timestamp 1668240031
transform -1 0 19964 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1019_
timestamp 1668240031
transform 1 0 17388 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1020_
timestamp 1668240031
transform -1 0 16376 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1021_
timestamp 1668240031
transform -1 0 15548 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1022_
timestamp 1668240031
transform 1 0 16836 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1023_
timestamp 1668240031
transform 1 0 12696 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1024_
timestamp 1668240031
transform -1 0 11224 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1025_
timestamp 1668240031
transform 1 0 10396 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1026_
timestamp 1668240031
transform -1 0 10120 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1027_
timestamp 1668240031
transform 1 0 14260 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1028_
timestamp 1668240031
transform -1 0 13800 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1029_
timestamp 1668240031
transform -1 0 16284 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1030_
timestamp 1668240031
transform 1 0 16652 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1031_
timestamp 1668240031
transform -1 0 16284 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1032_
timestamp 1668240031
transform -1 0 16560 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1033_
timestamp 1668240031
transform 1 0 12236 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1034_
timestamp 1668240031
transform -1 0 11868 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1035_
timestamp 1668240031
transform -1 0 12880 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1036_
timestamp 1668240031
transform 1 0 11684 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1037_
timestamp 1668240031
transform -1 0 11408 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1038_
timestamp 1668240031
transform 1 0 11684 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1039_
timestamp 1668240031
transform -1 0 11960 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1040_
timestamp 1668240031
transform 1 0 9108 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1041_
timestamp 1668240031
transform -1 0 8556 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1042_
timestamp 1668240031
transform 1 0 9108 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1043_
timestamp 1668240031
transform 1 0 7636 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1044_
timestamp 1668240031
transform 1 0 8464 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1045_
timestamp 1668240031
transform -1 0 8648 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1046_
timestamp 1668240031
transform 1 0 6716 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1047_
timestamp 1668240031
transform -1 0 6072 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1048_
timestamp 1668240031
transform 1 0 6532 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1049_
timestamp 1668240031
transform 1 0 6348 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1050_
timestamp 1668240031
transform 1 0 6532 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1051_
timestamp 1668240031
transform -1 0 5704 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1052_
timestamp 1668240031
transform 1 0 6348 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1053_
timestamp 1668240031
transform -1 0 6072 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1054_
timestamp 1668240031
transform 1 0 8740 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1055_
timestamp 1668240031
transform -1 0 8280 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1056_
timestamp 1668240031
transform -1 0 16468 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1057_
timestamp 1668240031
transform -1 0 13708 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1058_
timestamp 1668240031
transform 1 0 13432 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1059_
timestamp 1668240031
transform -1 0 12144 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1060_
timestamp 1668240031
transform 1 0 11684 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1061_
timestamp 1668240031
transform 1 0 9844 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1062_
timestamp 1668240031
transform 1 0 9936 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1063_
timestamp 1668240031
transform 1 0 7820 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1064_
timestamp 1668240031
transform -1 0 6256 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1065_
timestamp 1668240031
transform 1 0 7820 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1066_
timestamp 1668240031
transform 1 0 7728 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1067_
timestamp 1668240031
transform 1 0 9660 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1068_
timestamp 1668240031
transform -1 0 8648 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1069_
timestamp 1668240031
transform 1 0 11684 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1070_
timestamp 1668240031
transform -1 0 10764 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1071_
timestamp 1668240031
transform -1 0 13708 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1072_
timestamp 1668240031
transform 1 0 13340 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1073_
timestamp 1668240031
transform -1 0 13984 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1074_
timestamp 1668240031
transform -1 0 14168 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1075_
timestamp 1668240031
transform 1 0 14260 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1076_
timestamp 1668240031
transform -1 0 14536 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1077_
timestamp 1668240031
transform -1 0 16652 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1078_
timestamp 1668240031
transform 1 0 17204 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1079_
timestamp 1668240031
transform 1 0 14812 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1080_
timestamp 1668240031
transform -1 0 13800 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1081_
timestamp 1668240031
transform 1 0 17020 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1082_
timestamp 1668240031
transform -1 0 15732 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1083_
timestamp 1668240031
transform 1 0 19044 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1084_
timestamp 1668240031
transform -1 0 16376 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1085_
timestamp 1668240031
transform 1 0 20608 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1086_
timestamp 1668240031
transform -1 0 20884 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1087_
timestamp 1668240031
transform 1 0 20148 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1088_
timestamp 1668240031
transform -1 0 19964 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1089_
timestamp 1668240031
transform -1 0 20424 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1090_
timestamp 1668240031
transform 1 0 19964 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1091_
timestamp 1668240031
transform 1 0 19504 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1092_
timestamp 1668240031
transform -1 0 19320 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1093_
timestamp 1668240031
transform 1 0 18124 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1094_
timestamp 1668240031
transform -1 0 18308 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1095_
timestamp 1668240031
transform 1 0 16836 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1096_
timestamp 1668240031
transform 1 0 16100 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1097_
timestamp 1668240031
transform 1 0 14168 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1098_
timestamp 1668240031
transform 1 0 13524 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1099_
timestamp 1668240031
transform 1 0 12420 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1100_
timestamp 1668240031
transform 1 0 12696 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1101_
timestamp 1668240031
transform -1 0 11408 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1102_
timestamp 1668240031
transform 1 0 9568 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1103_
timestamp 1668240031
transform -1 0 9844 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1104_
timestamp 1668240031
transform 1 0 7820 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1105_
timestamp 1668240031
transform -1 0 6164 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1106_
timestamp 1668240031
transform 1 0 7820 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1107_
timestamp 1668240031
transform -1 0 6808 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1108_
timestamp 1668240031
transform 1 0 10396 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1109_
timestamp 1668240031
transform -1 0 9384 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1110_
timestamp 1668240031
transform 1 0 11776 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1111_
timestamp 1668240031
transform -1 0 11224 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1112_
timestamp 1668240031
transform 1 0 12604 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1113_
timestamp 1668240031
transform -1 0 11868 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1114_
timestamp 1668240031
transform 1 0 7820 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1115_
timestamp 1668240031
transform 1 0 7176 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1116_
timestamp 1668240031
transform 1 0 7820 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1117_
timestamp 1668240031
transform -1 0 6808 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1118_
timestamp 1668240031
transform 1 0 9568 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1119_
timestamp 1668240031
transform 1 0 9384 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1120_
timestamp 1668240031
transform -1 0 14812 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1121_
timestamp 1668240031
transform 1 0 12604 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1122_
timestamp 1668240031
transform -1 0 11224 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1123_
timestamp 1668240031
transform 1 0 14536 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1124_
timestamp 1668240031
transform 1 0 14444 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1125_
timestamp 1668240031
transform 1 0 15548 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1126_
timestamp 1668240031
transform -1 0 15180 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1127_
timestamp 1668240031
transform 1 0 16836 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1128_
timestamp 1668240031
transform 1 0 16836 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1129_
timestamp 1668240031
transform 1 0 19412 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1130_
timestamp 1668240031
transform 1 0 19412 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1131_
timestamp 1668240031
transform 1 0 19504 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1132_
timestamp 1668240031
transform -1 0 18952 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1133_
timestamp 1668240031
transform 1 0 16928 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1134_
timestamp 1668240031
transform 1 0 16100 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1135_
timestamp 1668240031
transform -1 0 21436 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1136_
timestamp 1668240031
transform -1 0 21160 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1137_
timestamp 1668240031
transform 1 0 19688 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1138_
timestamp 1668240031
transform -1 0 19872 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1139_
timestamp 1668240031
transform 1 0 19412 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1140_
timestamp 1668240031
transform -1 0 18308 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1141_
timestamp 1668240031
transform -1 0 26404 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1142_
timestamp 1668240031
transform -1 0 25392 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1143_
timestamp 1668240031
transform 1 0 25760 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1144_
timestamp 1668240031
transform 1 0 25484 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1145_
timestamp 1668240031
transform 1 0 25208 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1146_
timestamp 1668240031
transform -1 0 25392 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1147_
timestamp 1668240031
transform 1 0 26220 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1148_
timestamp 1668240031
transform 1 0 24564 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1149_
timestamp 1668240031
transform -1 0 24472 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1150_
timestamp 1668240031
transform -1 0 25300 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1151_
timestamp 1668240031
transform 1 0 25668 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1152_
timestamp 1668240031
transform 1 0 24564 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1153_
timestamp 1668240031
transform -1 0 24288 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1154_
timestamp 1668240031
transform -1 0 25484 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1155_
timestamp 1668240031
transform 1 0 25760 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1156_
timestamp 1668240031
transform -1 0 25392 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1157_
timestamp 1668240031
transform 1 0 25760 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1158_
timestamp 1668240031
transform -1 0 25208 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1159_
timestamp 1668240031
transform 1 0 25576 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1160_
timestamp 1668240031
transform -1 0 25852 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1161_
timestamp 1668240031
transform -1 0 26496 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1162_
timestamp 1668240031
transform -1 0 26128 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1163_
timestamp 1668240031
transform 1 0 24656 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1164_
timestamp 1668240031
transform -1 0 26680 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1165_
timestamp 1668240031
transform 1 0 27692 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1166_
timestamp 1668240031
transform -1 0 27140 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1167_
timestamp 1668240031
transform 1 0 27140 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1168_
timestamp 1668240031
transform -1 0 26588 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1169_
timestamp 1668240031
transform -1 0 26588 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1170_
timestamp 1668240031
transform -1 0 26404 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1171_
timestamp 1668240031
transform -1 0 26404 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1172_
timestamp 1668240031
transform -1 0 26588 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1173_
timestamp 1668240031
transform -1 0 26680 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1174_
timestamp 1668240031
transform 1 0 27140 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1175_
timestamp 1668240031
transform -1 0 26680 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1176_
timestamp 1668240031
transform -1 0 26312 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1177_
timestamp 1668240031
transform -1 0 27048 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1178_
timestamp 1668240031
transform -1 0 26036 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1179_
timestamp 1668240031
transform -1 0 26312 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1180_
timestamp 1668240031
transform 1 0 25392 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1181_
timestamp 1668240031
transform -1 0 24840 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1182_
timestamp 1668240031
transform -1 0 26220 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1183_
timestamp 1668240031
transform 1 0 28336 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1184_
timestamp 1668240031
transform 1 0 25760 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1185_
timestamp 1668240031
transform 1 0 27140 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1186_
timestamp 1668240031
transform -1 0 24104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1187_
timestamp 1668240031
transform 1 0 24564 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1188_
timestamp 1668240031
transform -1 0 24840 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1189_
timestamp 1668240031
transform 1 0 24196 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1190_
timestamp 1668240031
transform -1 0 24104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1191_
timestamp 1668240031
transform -1 0 27968 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1192_
timestamp 1668240031
transform 1 0 28796 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1193_
timestamp 1668240031
transform -1 0 28244 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1194_
timestamp 1668240031
transform 1 0 28888 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1195_
timestamp 1668240031
transform 1 0 29716 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1196_
timestamp 1668240031
transform 1 0 29716 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1197_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1668240031
transform 1 0 27784 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1198_
timestamp 1668240031
transform 1 0 27416 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1199_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1668240031
transform 1 0 30544 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1200_
timestamp 1668240031
transform 1 0 28060 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1201_
timestamp 1668240031
transform 1 0 28704 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1202_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1668240031
transform 1 0 29624 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1203_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1668240031
transform -1 0 30268 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1204_
timestamp 1668240031
transform 1 0 28428 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1205_
timestamp 1668240031
transform -1 0 28060 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__a21boi_1  _1206_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1668240031
transform 1 0 27600 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__o22ai_1  _1207_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1668240031
transform 1 0 28980 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _1208_
timestamp 1668240031
transform -1 0 28060 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1209_
timestamp 1668240031
transform 1 0 28152 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1210_
timestamp 1668240031
transform 1 0 27232 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1211_
timestamp 1668240031
transform -1 0 29624 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _1212_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1668240031
transform 1 0 27692 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1213_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1668240031
transform 1 0 27140 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1214_
timestamp 1668240031
transform 1 0 27968 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1215_
timestamp 1668240031
transform 1 0 27600 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1216_
timestamp 1668240031
transform -1 0 29072 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__a2111o_1  _1217_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1668240031
transform -1 0 28704 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__or2b_1  _1218_
timestamp 1668240031
transform -1 0 30268 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1219_
timestamp 1668240031
transform 1 0 26956 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1220_
timestamp 1668240031
transform -1 0 30268 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__o2111a_1  _1221_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1668240031
transform -1 0 28704 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _1222_
timestamp 1668240031
transform 1 0 28796 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _1223_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1668240031
transform 1 0 27784 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_1  _1224_
timestamp 1668240031
transform -1 0 29256 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__a41o_1  _1225_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1668240031
transform -1 0 28428 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1226_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1668240031
transform -1 0 28980 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1227_
timestamp 1668240031
transform -1 0 32568 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1228_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1668240031
transform -1 0 29900 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1229_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1668240031
transform -1 0 29256 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__nand3b_1  _1230_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1668240031
transform 1 0 29716 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1231_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1668240031
transform 1 0 31188 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1232_
timestamp 1668240031
transform -1 0 32568 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1233_
timestamp 1668240031
transform 1 0 32292 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1234_
timestamp 1668240031
transform -1 0 31832 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1235_
timestamp 1668240031
transform -1 0 30176 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1236_
timestamp 1668240031
transform 1 0 30544 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1237_
timestamp 1668240031
transform -1 0 29992 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1238_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1668240031
transform 1 0 32292 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1239_
timestamp 1668240031
transform -1 0 32476 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1240_
timestamp 1668240031
transform 1 0 31004 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1241_
timestamp 1668240031
transform 1 0 32292 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1242_
timestamp 1668240031
transform 1 0 32200 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1243_
timestamp 1668240031
transform -1 0 33580 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1244_
timestamp 1668240031
transform 1 0 33304 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1245_
timestamp 1668240031
transform 1 0 30728 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1246_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1668240031
transform -1 0 30268 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_2  _1247_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1668240031
transform -1 0 31280 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1248_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1668240031
transform 1 0 32200 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1249_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1668240031
transform -1 0 33396 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1250_
timestamp 1668240031
transform 1 0 32200 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1251_
timestamp 1668240031
transform 1 0 32292 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1252_
timestamp 1668240031
transform 1 0 33580 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1253_
timestamp 1668240031
transform 1 0 32752 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1254_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1668240031
transform -1 0 33856 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1255_
timestamp 1668240031
transform 1 0 32292 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1256_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1668240031
transform 1 0 29348 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1257_
timestamp 1668240031
transform -1 0 29256 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1258_
timestamp 1668240031
transform 1 0 28612 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1259_
timestamp 1668240031
transform 1 0 28428 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1260_
timestamp 1668240031
transform -1 0 34040 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1261_
timestamp 1668240031
transform -1 0 31832 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1262_
timestamp 1668240031
transform 1 0 30176 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1263_
timestamp 1668240031
transform 1 0 29716 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1264_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1668240031
transform -1 0 29900 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1265_
timestamp 1668240031
transform -1 0 32752 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1266_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1668240031
transform -1 0 29256 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1267_
timestamp 1668240031
transform -1 0 29072 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1268_
timestamp 1668240031
transform -1 0 29624 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _1269_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1668240031
transform 1 0 28244 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1270_
timestamp 1668240031
transform 1 0 28520 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1271_
timestamp 1668240031
transform -1 0 30084 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1272_
timestamp 1668240031
transform 1 0 28152 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1273_
timestamp 1668240031
transform -1 0 34132 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1274_
timestamp 1668240031
transform 1 0 27784 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1275_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1668240031
transform 1 0 27140 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1276_
timestamp 1668240031
transform 1 0 28336 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1277_
timestamp 1668240031
transform 1 0 29716 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1278_
timestamp 1668240031
transform 1 0 28520 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1279_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1668240031
transform 1 0 28152 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1280_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1668240031
transform 1 0 28428 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_1  _1281_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1668240031
transform 1 0 29716 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1282_
timestamp 1668240031
transform 1 0 30544 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1283_
timestamp 1668240031
transform 1 0 27416 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1284_
timestamp 1668240031
transform -1 0 29348 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1285_
timestamp 1668240031
transform -1 0 29992 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1286_
timestamp 1668240031
transform -1 0 27416 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1287_
timestamp 1668240031
transform 1 0 31464 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1288_
timestamp 1668240031
transform -1 0 30912 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1289_
timestamp 1668240031
transform 1 0 27232 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1290_
timestamp 1668240031
transform 1 0 27324 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1291_
timestamp 1668240031
transform 1 0 27692 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _1292_
timestamp 1668240031
transform -1 0 29072 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1293_
timestamp 1668240031
transform 1 0 28336 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1294_
timestamp 1668240031
transform -1 0 30912 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1295_
timestamp 1668240031
transform 1 0 28336 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1296_
timestamp 1668240031
transform 1 0 27692 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1297_
timestamp 1668240031
transform -1 0 30360 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1298_
timestamp 1668240031
transform -1 0 28888 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _1299_
timestamp 1668240031
transform -1 0 29348 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1300_
timestamp 1668240031
transform 1 0 28244 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _1301_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1668240031
transform -1 0 29256 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _1302_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1668240031
transform 1 0 29532 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1303_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1668240031
transform 1 0 29716 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1304_
timestamp 1668240031
transform 1 0 31096 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1305_
timestamp 1668240031
transform 1 0 31372 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1306_
timestamp 1668240031
transform -1 0 32844 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1307_
timestamp 1668240031
transform 1 0 28520 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _1308_
timestamp 1668240031
transform 1 0 28428 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1309_
timestamp 1668240031
transform 1 0 28704 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _1310_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1668240031
transform 1 0 30360 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _1311_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1668240031
transform 1 0 29348 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_4  _1312_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1668240031
transform 1 0 29716 0 1 25024
box -38 -48 1326 592
use sky130_fd_sc_hd__mux2_1  _1313_
timestamp 1668240031
transform -1 0 30268 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1314_
timestamp 1668240031
transform 1 0 31280 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1315_
timestamp 1668240031
transform 1 0 29716 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1316_
timestamp 1668240031
transform -1 0 30912 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1317_
timestamp 1668240031
transform 1 0 30636 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1318_
timestamp 1668240031
transform -1 0 34040 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1319_
timestamp 1668240031
transform -1 0 35328 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1320_
timestamp 1668240031
transform -1 0 33028 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1321_
timestamp 1668240031
transform 1 0 33580 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1322_
timestamp 1668240031
transform 1 0 34868 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1323_
timestamp 1668240031
transform -1 0 35236 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1324_
timestamp 1668240031
transform 1 0 33304 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1325_
timestamp 1668240031
transform -1 0 34224 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1326_
timestamp 1668240031
transform 1 0 34316 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1327_
timestamp 1668240031
transform 1 0 34040 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _1328_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1668240031
transform -1 0 34224 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _1329_
timestamp 1668240031
transform 1 0 33304 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1330_
timestamp 1668240031
transform 1 0 34868 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1331_
timestamp 1668240031
transform -1 0 34684 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1332_
timestamp 1668240031
transform 1 0 33212 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1333_
timestamp 1668240031
transform -1 0 35328 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1334_
timestamp 1668240031
transform -1 0 35236 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1335_
timestamp 1668240031
transform -1 0 35972 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1336_
timestamp 1668240031
transform -1 0 36708 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _1337_
timestamp 1668240031
transform -1 0 33856 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1338_
timestamp 1668240031
transform 1 0 33764 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1339_
timestamp 1668240031
transform -1 0 35052 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1340_
timestamp 1668240031
transform -1 0 35972 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1341_
timestamp 1668240031
transform 1 0 33304 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1342_
timestamp 1668240031
transform -1 0 35696 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1343_
timestamp 1668240031
transform 1 0 35512 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1344_
timestamp 1668240031
transform -1 0 34224 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1345_
timestamp 1668240031
transform 1 0 34868 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1346_
timestamp 1668240031
transform 1 0 30176 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1347_
timestamp 1668240031
transform -1 0 31188 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1348_
timestamp 1668240031
transform -1 0 31832 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1349_
timestamp 1668240031
transform -1 0 36064 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _1350_
timestamp 1668240031
transform -1 0 14812 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1351_
timestamp 1668240031
transform 1 0 28612 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1352_
timestamp 1668240031
transform 1 0 30360 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1353_
timestamp 1668240031
transform -1 0 30544 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1354_
timestamp 1668240031
transform 1 0 31188 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1355_
timestamp 1668240031
transform 1 0 28428 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1356_
timestamp 1668240031
transform 1 0 27140 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1357_
timestamp 1668240031
transform 1 0 27140 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1358_
timestamp 1668240031
transform -1 0 28336 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1359_
timestamp 1668240031
transform -1 0 30544 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1360_
timestamp 1668240031
transform 1 0 30912 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1361_
timestamp 1668240031
transform 1 0 30268 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1362_
timestamp 1668240031
transform -1 0 30544 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1363_
timestamp 1668240031
transform 1 0 33948 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1364_
timestamp 1668240031
transform 1 0 31556 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  _1365_
timestamp 1668240031
transform -1 0 17848 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1366_
timestamp 1668240031
transform -1 0 31832 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1367_
timestamp 1668240031
transform -1 0 31740 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1368_
timestamp 1668240031
transform 1 0 32752 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1369_
timestamp 1668240031
transform -1 0 31832 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1370_
timestamp 1668240031
transform 1 0 33304 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1371_
timestamp 1668240031
transform 1 0 32108 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1372_
timestamp 1668240031
transform 1 0 31372 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1373_
timestamp 1668240031
transform 1 0 31464 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1374_
timestamp 1668240031
transform 1 0 33488 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1375_
timestamp 1668240031
transform -1 0 33120 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1376_
timestamp 1668240031
transform 1 0 34868 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1377_
timestamp 1668240031
transform -1 0 32936 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1378_
timestamp 1668240031
transform 1 0 32292 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1379_
timestamp 1668240031
transform 1 0 31924 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1380_
timestamp 1668240031
transform 1 0 29164 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1381_
timestamp 1668240031
transform 1 0 28152 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1382_
timestamp 1668240031
transform 1 0 27508 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1383_
timestamp 1668240031
transform -1 0 23736 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1384_
timestamp 1668240031
transform 1 0 24196 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1385_
timestamp 1668240031
transform 1 0 22448 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1386_
timestamp 1668240031
transform -1 0 22080 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1387_
timestamp 1668240031
transform 1 0 22448 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1388_
timestamp 1668240031
transform 1 0 20332 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1389_
timestamp 1668240031
transform 1 0 19780 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1390_
timestamp 1668240031
transform 1 0 18124 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1391_
timestamp 1668240031
transform 1 0 18032 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1392_
timestamp 1668240031
transform 1 0 17480 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1393_
timestamp 1668240031
transform 1 0 16284 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1394_
timestamp 1668240031
transform 1 0 15916 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1395_
timestamp 1668240031
transform 1 0 15456 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1396_
timestamp 1668240031
transform 1 0 13340 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _1397_
timestamp 1668240031
transform 1 0 14260 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1398_
timestamp 1668240031
transform 1 0 10948 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1399_
timestamp 1668240031
transform -1 0 10580 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1400_
timestamp 1668240031
transform -1 0 12972 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1401_
timestamp 1668240031
transform 1 0 12144 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1402_
timestamp 1668240031
transform 1 0 11776 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1403_
timestamp 1668240031
transform -1 0 13432 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1404_
timestamp 1668240031
transform 1 0 12604 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1405_
timestamp 1668240031
transform 1 0 12144 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1406_
timestamp 1668240031
transform 1 0 14260 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1407_
timestamp 1668240031
transform -1 0 15088 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1408_
timestamp 1668240031
transform 1 0 15732 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1409_
timestamp 1668240031
transform 1 0 15088 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1410_
timestamp 1668240031
transform 1 0 14076 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1411_
timestamp 1668240031
transform -1 0 13708 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1412_
timestamp 1668240031
transform 1 0 13892 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1413_
timestamp 1668240031
transform 1 0 12052 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1414_
timestamp 1668240031
transform -1 0 11224 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1415_
timestamp 1668240031
transform -1 0 13616 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1416_
timestamp 1668240031
transform 1 0 12328 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1417_
timestamp 1668240031
transform -1 0 11224 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1418_
timestamp 1668240031
transform 1 0 10672 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1419_
timestamp 1668240031
transform 1 0 10488 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1420_
timestamp 1668240031
transform 1 0 10396 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1421_
timestamp 1668240031
transform -1 0 10764 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1422_
timestamp 1668240031
transform 1 0 9292 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1423_
timestamp 1668240031
transform 1 0 9108 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1424_
timestamp 1668240031
transform -1 0 8648 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1425_
timestamp 1668240031
transform 1 0 9108 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1426_
timestamp 1668240031
transform 1 0 9016 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1427_
timestamp 1668240031
transform -1 0 8648 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1428_
timestamp 1668240031
transform 1 0 9660 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  _1429_
timestamp 1668240031
transform -1 0 13800 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1430_
timestamp 1668240031
transform -1 0 10304 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1431_
timestamp 1668240031
transform 1 0 11316 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1432_
timestamp 1668240031
transform 1 0 7820 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1433_
timestamp 1668240031
transform -1 0 7452 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1434_
timestamp 1668240031
transform -1 0 8188 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1435_
timestamp 1668240031
transform 1 0 6992 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1436_
timestamp 1668240031
transform 1 0 6532 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1437_
timestamp 1668240031
transform -1 0 6440 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1438_
timestamp 1668240031
transform 1 0 6992 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1439_
timestamp 1668240031
transform 1 0 6624 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1440_
timestamp 1668240031
transform -1 0 6072 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1441_
timestamp 1668240031
transform 1 0 7544 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1442_
timestamp 1668240031
transform 1 0 6440 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1443_
timestamp 1668240031
transform -1 0 6072 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1444_
timestamp 1668240031
transform 1 0 9936 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1445_
timestamp 1668240031
transform 1 0 8556 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1446_
timestamp 1668240031
transform -1 0 8188 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1447_
timestamp 1668240031
transform -1 0 13892 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1448_
timestamp 1668240031
transform 1 0 12236 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1449_
timestamp 1668240031
transform 1 0 11684 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1450_
timestamp 1668240031
transform -1 0 11224 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1451_
timestamp 1668240031
transform 1 0 11684 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1452_
timestamp 1668240031
transform 1 0 10120 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1453_
timestamp 1668240031
transform -1 0 9016 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1454_
timestamp 1668240031
transform 1 0 11040 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1455_
timestamp 1668240031
transform 1 0 10212 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1456_
timestamp 1668240031
transform 1 0 8372 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1457_
timestamp 1668240031
transform 1 0 9108 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1458_
timestamp 1668240031
transform 1 0 8004 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1459_
timestamp 1668240031
transform 1 0 7360 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1460_
timestamp 1668240031
transform 1 0 9108 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _1461_
timestamp 1668240031
transform -1 0 14812 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1462_
timestamp 1668240031
transform -1 0 7452 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1463_
timestamp 1668240031
transform 1 0 7268 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1464_
timestamp 1668240031
transform 1 0 9292 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1465_
timestamp 1668240031
transform 1 0 9200 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1466_
timestamp 1668240031
transform -1 0 9568 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1467_
timestamp 1668240031
transform -1 0 11224 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1468_
timestamp 1668240031
transform 1 0 10396 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1469_
timestamp 1668240031
transform -1 0 10856 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1470_
timestamp 1668240031
transform -1 0 12604 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1471_
timestamp 1668240031
transform 1 0 12696 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1472_
timestamp 1668240031
transform -1 0 11592 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1473_
timestamp 1668240031
transform 1 0 12512 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1474_
timestamp 1668240031
transform 1 0 12052 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1475_
timestamp 1668240031
transform -1 0 11684 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1476_
timestamp 1668240031
transform -1 0 13800 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1477_
timestamp 1668240031
transform 1 0 12972 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1478_
timestamp 1668240031
transform -1 0 12604 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1479_
timestamp 1668240031
transform 1 0 15364 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1480_
timestamp 1668240031
transform 1 0 14904 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1481_
timestamp 1668240031
transform -1 0 15548 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1482_
timestamp 1668240031
transform 1 0 15180 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1483_
timestamp 1668240031
transform -1 0 17664 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1484_
timestamp 1668240031
transform 1 0 16836 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1485_
timestamp 1668240031
transform -1 0 17204 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1486_
timestamp 1668240031
transform -1 0 18952 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1487_
timestamp 1668240031
transform -1 0 19320 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1488_
timestamp 1668240031
transform -1 0 19136 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1489_
timestamp 1668240031
transform 1 0 20332 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1490_
timestamp 1668240031
transform -1 0 20792 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1491_
timestamp 1668240031
transform 1 0 21160 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1492_
timestamp 1668240031
transform 1 0 20424 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _1493_
timestamp 1668240031
transform 1 0 14812 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1494_
timestamp 1668240031
transform -1 0 18952 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1495_
timestamp 1668240031
transform -1 0 19688 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1496_
timestamp 1668240031
transform 1 0 19504 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1497_
timestamp 1668240031
transform 1 0 18676 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1498_
timestamp 1668240031
transform 1 0 18124 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1499_
timestamp 1668240031
transform 1 0 19412 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1500_
timestamp 1668240031
transform -1 0 18952 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1501_
timestamp 1668240031
transform 1 0 20608 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1502_
timestamp 1668240031
transform -1 0 18952 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1503_
timestamp 1668240031
transform -1 0 18952 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1504_
timestamp 1668240031
transform 1 0 20056 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1505_
timestamp 1668240031
transform 1 0 16836 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1506_
timestamp 1668240031
transform 1 0 15732 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1507_
timestamp 1668240031
transform 1 0 15272 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1508_
timestamp 1668240031
transform 1 0 15364 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1509_
timestamp 1668240031
transform 1 0 14260 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1510_
timestamp 1668240031
transform -1 0 10580 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1511_
timestamp 1668240031
transform -1 0 13800 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1512_
timestamp 1668240031
transform 1 0 12328 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1513_
timestamp 1668240031
transform -1 0 11776 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1514_
timestamp 1668240031
transform 1 0 11684 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1515_
timestamp 1668240031
transform 1 0 11684 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1516_
timestamp 1668240031
transform 1 0 7820 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1517_
timestamp 1668240031
transform 1 0 7728 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1518_
timestamp 1668240031
transform 1 0 9108 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1519_
timestamp 1668240031
transform 1 0 7728 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1520_
timestamp 1668240031
transform 1 0 6992 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1521_
timestamp 1668240031
transform 1 0 8004 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1522_
timestamp 1668240031
transform 1 0 6808 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1523_
timestamp 1668240031
transform -1 0 7268 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1524_
timestamp 1668240031
transform -1 0 10028 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _1525_
timestamp 1668240031
transform 1 0 14352 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1526_
timestamp 1668240031
transform 1 0 9752 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1527_
timestamp 1668240031
transform -1 0 7452 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1528_
timestamp 1668240031
transform 1 0 11684 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1529_
timestamp 1668240031
transform 1 0 10396 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1530_
timestamp 1668240031
transform -1 0 8740 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1531_
timestamp 1668240031
transform -1 0 12420 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1532_
timestamp 1668240031
transform 1 0 11684 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1533_
timestamp 1668240031
transform -1 0 10580 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1534_
timestamp 1668240031
transform 1 0 9568 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1535_
timestamp 1668240031
transform 1 0 9108 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1536_
timestamp 1668240031
transform -1 0 7452 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1537_
timestamp 1668240031
transform 1 0 9108 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1538_
timestamp 1668240031
transform 1 0 8464 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1539_
timestamp 1668240031
transform -1 0 7452 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1540_
timestamp 1668240031
transform 1 0 11684 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1541_
timestamp 1668240031
transform -1 0 11224 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1542_
timestamp 1668240031
transform -1 0 11040 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1543_
timestamp 1668240031
transform -1 0 19964 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1544_
timestamp 1668240031
transform 1 0 12972 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1545_
timestamp 1668240031
transform -1 0 13708 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1546_
timestamp 1668240031
transform 1 0 16100 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1547_
timestamp 1668240031
transform -1 0 15640 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1548_
timestamp 1668240031
transform 1 0 14904 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1549_
timestamp 1668240031
transform -1 0 13800 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1550_
timestamp 1668240031
transform 1 0 15548 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1551_
timestamp 1668240031
transform 1 0 14628 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1552_
timestamp 1668240031
transform -1 0 14536 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1553_
timestamp 1668240031
transform 1 0 15548 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1554_
timestamp 1668240031
transform 1 0 14720 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1555_
timestamp 1668240031
transform -1 0 11960 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1556_
timestamp 1668240031
transform 1 0 18676 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _1557_
timestamp 1668240031
transform -1 0 20884 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1558_
timestamp 1668240031
transform 1 0 17480 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1559_
timestamp 1668240031
transform -1 0 17112 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1560_
timestamp 1668240031
transform 1 0 19136 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1561_
timestamp 1668240031
transform 1 0 18124 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1562_
timestamp 1668240031
transform -1 0 17664 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1563_
timestamp 1668240031
transform 1 0 18032 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1564_
timestamp 1668240031
transform 1 0 17480 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1565_
timestamp 1668240031
transform -1 0 16376 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1566_
timestamp 1668240031
transform 1 0 18124 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1567_
timestamp 1668240031
transform 1 0 17756 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1568_
timestamp 1668240031
transform 1 0 17112 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1569_
timestamp 1668240031
transform 1 0 19412 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1570_
timestamp 1668240031
transform -1 0 18952 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1571_
timestamp 1668240031
transform 1 0 20332 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1572_
timestamp 1668240031
transform -1 0 20516 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1573_
timestamp 1668240031
transform -1 0 20608 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1574_
timestamp 1668240031
transform 1 0 20976 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1575_
timestamp 1668240031
transform 1 0 22908 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1576_
timestamp 1668240031
transform 1 0 23460 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1577_
timestamp 1668240031
transform 1 0 23000 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1578_
timestamp 1668240031
transform 1 0 22540 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1579_
timestamp 1668240031
transform 1 0 24288 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1580_
timestamp 1668240031
transform -1 0 24104 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1581_
timestamp 1668240031
transform 1 0 24564 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1582_
timestamp 1668240031
transform 1 0 25760 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1583_
timestamp 1668240031
transform 1 0 23276 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1584_
timestamp 1668240031
transform 1 0 22724 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1585_
timestamp 1668240031
transform 1 0 24380 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1586_
timestamp 1668240031
transform 1 0 22816 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1587_
timestamp 1668240031
transform 1 0 22632 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1588_
timestamp 1668240031
transform 1 0 23184 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _1589_
timestamp 1668240031
transform 1 0 22724 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1590_
timestamp 1668240031
transform 1 0 22908 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1591_
timestamp 1668240031
transform 1 0 21988 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1592_
timestamp 1668240031
transform 1 0 23276 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1593_
timestamp 1668240031
transform -1 0 23276 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1594_
timestamp 1668240031
transform 1 0 23368 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1595_
timestamp 1668240031
transform 1 0 23460 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1596_
timestamp 1668240031
transform 1 0 23092 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1597_
timestamp 1668240031
transform 1 0 21252 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1598_
timestamp 1668240031
transform 1 0 23552 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1599_
timestamp 1668240031
transform 1 0 22356 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1600_
timestamp 1668240031
transform 1 0 20884 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1601_
timestamp 1668240031
transform 1 0 23184 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1602_
timestamp 1668240031
transform 1 0 22172 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1603_
timestamp 1668240031
transform 1 0 21988 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1604_
timestamp 1668240031
transform 1 0 23828 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1605_
timestamp 1668240031
transform -1 0 24012 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1606_
timestamp 1668240031
transform 1 0 24564 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1607_
timestamp 1668240031
transform 1 0 24564 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1608_
timestamp 1668240031
transform 1 0 24472 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1609_
timestamp 1668240031
transform 1 0 23276 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1610_
timestamp 1668240031
transform 1 0 22448 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1611_
timestamp 1668240031
transform 1 0 25668 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1612_
timestamp 1668240031
transform -1 0 25392 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1613_
timestamp 1668240031
transform 1 0 26404 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1614_
timestamp 1668240031
transform 1 0 25116 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1615_
timestamp 1668240031
transform 1 0 24012 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1616_
timestamp 1668240031
transform 1 0 22908 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1617_
timestamp 1668240031
transform 1 0 25024 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1618_
timestamp 1668240031
transform 1 0 24932 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1619_
timestamp 1668240031
transform 1 0 23828 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1620_
timestamp 1668240031
transform 1 0 25208 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _1621_
timestamp 1668240031
transform -1 0 25116 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1622_
timestamp 1668240031
transform 1 0 24564 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1623_
timestamp 1668240031
transform 1 0 24564 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1624_
timestamp 1668240031
transform 1 0 25208 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1625_
timestamp 1668240031
transform 1 0 23276 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1626_
timestamp 1668240031
transform 1 0 22356 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1627_
timestamp 1668240031
transform 1 0 25760 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1628_
timestamp 1668240031
transform 1 0 24564 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1629_
timestamp 1668240031
transform -1 0 24104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1630_
timestamp 1668240031
transform 1 0 24840 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1631_
timestamp 1668240031
transform 1 0 23184 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1632_
timestamp 1668240031
transform 1 0 22540 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1633_
timestamp 1668240031
transform 1 0 24196 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1634_
timestamp 1668240031
transform 1 0 23000 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1635_
timestamp 1668240031
transform -1 0 22356 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1636_
timestamp 1668240031
transform 1 0 24196 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1637_
timestamp 1668240031
transform 1 0 23000 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1638_
timestamp 1668240031
transform 1 0 22172 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1639_
timestamp 1668240031
transform 1 0 23276 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1640_
timestamp 1668240031
transform -1 0 22908 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1641_
timestamp 1668240031
transform 1 0 23368 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1642_
timestamp 1668240031
transform 1 0 23184 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1643_
timestamp 1668240031
transform 1 0 22448 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1644_
timestamp 1668240031
transform 1 0 21712 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1645_
timestamp 1668240031
transform 1 0 24380 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1646_
timestamp 1668240031
transform 1 0 23276 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1647_
timestamp 1668240031
transform 1 0 22264 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1648_
timestamp 1668240031
transform -1 0 25392 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1649_
timestamp 1668240031
transform 1 0 25392 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1650_
timestamp 1668240031
transform 1 0 22540 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1651_
timestamp 1668240031
transform 1 0 26220 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1652_
timestamp 1668240031
transform 1 0 25484 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1653_
timestamp 1668240031
transform 1 0 24748 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1654_
timestamp 1668240031
transform 1 0 28336 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1655_
timestamp 1668240031
transform 1 0 27140 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1656_
timestamp 1668240031
transform 1 0 25300 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1657_
timestamp 1668240031
transform -1 0 34408 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1658_
timestamp 1668240031
transform -1 0 34776 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1659_
timestamp 1668240031
transform -1 0 34408 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1660_
timestamp 1668240031
transform -1 0 34684 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1661_
timestamp 1668240031
transform -1 0 33120 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1662_
timestamp 1668240031
transform -1 0 33856 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1663_
timestamp 1668240031
transform 1 0 14444 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1664_
timestamp 1668240031
transform -1 0 13524 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1665_
timestamp 1668240031
transform 1 0 15456 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1666_
timestamp 1668240031
transform 1 0 14352 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1667_
timestamp 1668240031
transform 1 0 16744 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1668_
timestamp 1668240031
transform -1 0 16376 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1669_
timestamp 1668240031
transform 1 0 19412 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1670_
timestamp 1668240031
transform -1 0 16376 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1671_
timestamp 1668240031
transform 1 0 20608 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1672_
timestamp 1668240031
transform -1 0 16376 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1673_
timestamp 1668240031
transform 1 0 20976 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1674_
timestamp 1668240031
transform -1 0 15272 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1675_
timestamp 1668240031
transform 1 0 21988 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1676_
timestamp 1668240031
transform -1 0 16376 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1677_
timestamp 1668240031
transform 1 0 21804 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1678_
timestamp 1668240031
transform -1 0 17112 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1679_
timestamp 1668240031
transform 1 0 19228 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1680_
timestamp 1668240031
transform -1 0 18860 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1681_
timestamp 1668240031
transform 1 0 16836 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1682_
timestamp 1668240031
transform -1 0 15916 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1683_
timestamp 1668240031
transform 1 0 13892 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1684_
timestamp 1668240031
transform 1 0 12880 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1685_
timestamp 1668240031
transform 1 0 12420 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1686_
timestamp 1668240031
transform 1 0 5060 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1687_
timestamp 1668240031
transform 1 0 9752 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1688_
timestamp 1668240031
transform 1 0 8096 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1689_
timestamp 1668240031
transform 1 0 10304 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1690_
timestamp 1668240031
transform 1 0 10120 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1691_
timestamp 1668240031
transform -1 0 10856 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1692_
timestamp 1668240031
transform -1 0 10580 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1693_
timestamp 1668240031
transform -1 0 15088 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1694_
timestamp 1668240031
transform -1 0 15824 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1695_
timestamp 1668240031
transform -1 0 15088 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1696_
timestamp 1668240031
transform -1 0 15364 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1697_
timestamp 1668240031
transform 1 0 12788 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1698_
timestamp 1668240031
transform -1 0 12052 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1699_
timestamp 1668240031
transform 1 0 30452 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1700_
timestamp 1668240031
transform -1 0 31280 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1701_
timestamp 1668240031
transform -1 0 31464 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1702_
timestamp 1668240031
transform 1 0 32936 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1703_
timestamp 1668240031
transform 1 0 30084 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1704_
timestamp 1668240031
transform -1 0 31464 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1705_
timestamp 1668240031
transform 1 0 32292 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1706_
timestamp 1668240031
transform 1 0 29716 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1707_
timestamp 1668240031
transform 1 0 29808 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1708_
timestamp 1668240031
transform -1 0 31096 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1709_
timestamp 1668240031
transform -1 0 31740 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1710_
timestamp 1668240031
transform 1 0 30636 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1711_
timestamp 1668240031
transform -1 0 30912 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1712_
timestamp 1668240031
transform -1 0 31740 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1713_
timestamp 1668240031
transform 1 0 29716 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1714_
timestamp 1668240031
transform 1 0 29716 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1715_
timestamp 1668240031
transform 1 0 28888 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1716_
timestamp 1668240031
transform -1 0 31464 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1717_
timestamp 1668240031
transform 1 0 29624 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1718_
timestamp 1668240031
transform 1 0 33396 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1719_
timestamp 1668240031
transform 1 0 34868 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1720_
timestamp 1668240031
transform -1 0 35236 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1721_
timestamp 1668240031
transform 1 0 35604 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1722_
timestamp 1668240031
transform 1 0 34500 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1723_
timestamp 1668240031
transform 1 0 35328 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1724_
timestamp 1668240031
transform -1 0 34316 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1725_
timestamp 1668240031
transform -1 0 36340 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1726_
timestamp 1668240031
transform 1 0 35052 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1727_
timestamp 1668240031
transform -1 0 32752 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1728_
timestamp 1668240031
transform 1 0 32384 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1729_
timestamp 1668240031
transform -1 0 32476 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1730_
timestamp 1668240031
transform 1 0 30728 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1731_
timestamp 1668240031
transform 1 0 31280 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1732_
timestamp 1668240031
transform -1 0 30912 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1733_
timestamp 1668240031
transform 1 0 29716 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1734_
timestamp 1668240031
transform -1 0 31188 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1735_
timestamp 1668240031
transform 1 0 32292 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1736_
timestamp 1668240031
transform -1 0 30084 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1737_
timestamp 1668240031
transform 1 0 30452 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__buf_4  _1738_
timestamp 1668240031
transform -1 0 22908 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1739_
timestamp 1668240031
transform 1 0 18400 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _1740_
timestamp 1668240031
transform -1 0 22172 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1741_
timestamp 1668240031
transform 1 0 26036 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1742_
timestamp 1668240031
transform 1 0 25392 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1743_
timestamp 1668240031
transform -1 0 23920 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1744_
timestamp 1668240031
transform 1 0 22908 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1745_
timestamp 1668240031
transform 1 0 22080 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1746_
timestamp 1668240031
transform -1 0 21528 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1747_
timestamp 1668240031
transform 1 0 22540 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1748_
timestamp 1668240031
transform 1 0 21896 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1749_
timestamp 1668240031
transform 1 0 22816 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1750_
timestamp 1668240031
transform 1 0 24196 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1751_
timestamp 1668240031
transform 1 0 23000 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1752_
timestamp 1668240031
transform -1 0 24472 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1753_
timestamp 1668240031
transform -1 0 24840 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1754_
timestamp 1668240031
transform 1 0 23552 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1755_
timestamp 1668240031
transform 1 0 23184 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1756_
timestamp 1668240031
transform 1 0 25760 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1757_
timestamp 1668240031
transform -1 0 23828 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1758_
timestamp 1668240031
transform -1 0 25484 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1759_
timestamp 1668240031
transform -1 0 22264 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1760_
timestamp 1668240031
transform -1 0 23644 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1761_
timestamp 1668240031
transform -1 0 21528 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1762_
timestamp 1668240031
transform -1 0 18952 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1763_
timestamp 1668240031
transform 1 0 21252 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1764_
timestamp 1668240031
transform 1 0 21252 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1765_
timestamp 1668240031
transform 1 0 22172 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1766_
timestamp 1668240031
transform 1 0 25576 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1767_
timestamp 1668240031
transform 1 0 23644 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1768_
timestamp 1668240031
transform 1 0 23000 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1769_
timestamp 1668240031
transform -1 0 22264 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1770_
timestamp 1668240031
transform -1 0 19320 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1771_
timestamp 1668240031
transform -1 0 17756 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1772_
timestamp 1668240031
transform -1 0 18952 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1773_
timestamp 1668240031
transform -1 0 18584 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1774_
timestamp 1668240031
transform 1 0 17388 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1775_
timestamp 1668240031
transform 1 0 18032 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1776_
timestamp 1668240031
transform 1 0 13340 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1777_
timestamp 1668240031
transform 1 0 10948 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1778_
timestamp 1668240031
transform -1 0 15732 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1779_
timestamp 1668240031
transform 1 0 12236 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1780_
timestamp 1668240031
transform -1 0 12144 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1781_
timestamp 1668240031
transform -1 0 9292 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1782_
timestamp 1668240031
transform -1 0 8096 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1783_
timestamp 1668240031
transform 1 0 10948 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1784_
timestamp 1668240031
transform 1 0 17020 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1785_
timestamp 1668240031
transform 1 0 10304 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1786_
timestamp 1668240031
transform 1 0 9200 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1787_
timestamp 1668240031
transform -1 0 9384 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1788_
timestamp 1668240031
transform -1 0 7452 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1789_
timestamp 1668240031
transform 1 0 8372 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1790_
timestamp 1668240031
transform 1 0 8740 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1791_
timestamp 1668240031
transform -1 0 13800 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1792_
timestamp 1668240031
transform 1 0 15456 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1793_
timestamp 1668240031
transform -1 0 19688 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1794_
timestamp 1668240031
transform 1 0 21252 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1795_
timestamp 1668240031
transform 1 0 17296 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1796_
timestamp 1668240031
transform 1 0 18492 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1797_
timestamp 1668240031
transform -1 0 19412 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1798_
timestamp 1668240031
transform 1 0 20240 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1799_
timestamp 1668240031
transform 1 0 19596 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1800_
timestamp 1668240031
transform -1 0 18216 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1801_
timestamp 1668240031
transform 1 0 15548 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1802_
timestamp 1668240031
transform 1 0 12880 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1803_
timestamp 1668240031
transform 1 0 12328 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1804_
timestamp 1668240031
transform -1 0 12144 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1805_
timestamp 1668240031
transform -1 0 12236 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1806_
timestamp 1668240031
transform 1 0 27140 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _1807_
timestamp 1668240031
transform -1 0 14812 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1808_
timestamp 1668240031
transform 1 0 9936 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1809_
timestamp 1668240031
transform -1 0 8188 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1810_
timestamp 1668240031
transform 1 0 7820 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1811_
timestamp 1668240031
transform -1 0 9384 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1812_
timestamp 1668240031
transform 1 0 9476 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1813_
timestamp 1668240031
transform 1 0 11592 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1814_
timestamp 1668240031
transform 1 0 10120 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1815_
timestamp 1668240031
transform 1 0 5796 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1816_
timestamp 1668240031
transform -1 0 5888 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1817_
timestamp 1668240031
transform 1 0 6532 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1818_
timestamp 1668240031
transform 1 0 13432 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1819_
timestamp 1668240031
transform -1 0 9384 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1820_
timestamp 1668240031
transform -1 0 10856 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1821_
timestamp 1668240031
transform 1 0 9476 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1822_
timestamp 1668240031
transform -1 0 8648 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1823_
timestamp 1668240031
transform 1 0 14260 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1824_
timestamp 1668240031
transform 1 0 10488 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1825_
timestamp 1668240031
transform 1 0 11960 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1826_
timestamp 1668240031
transform 1 0 13524 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1827_
timestamp 1668240031
transform 1 0 14260 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1828_
timestamp 1668240031
transform 1 0 12788 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1829_
timestamp 1668240031
transform -1 0 17940 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1830_
timestamp 1668240031
transform 1 0 10948 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1831_
timestamp 1668240031
transform -1 0 10580 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1832_
timestamp 1668240031
transform -1 0 16284 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1833_
timestamp 1668240031
transform -1 0 18492 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1834_
timestamp 1668240031
transform -1 0 20700 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1835_
timestamp 1668240031
transform -1 0 23920 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1836_
timestamp 1668240031
transform 1 0 27968 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1837_
timestamp 1668240031
transform -1 0 32844 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1838_
timestamp 1668240031
transform 1 0 33304 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1839_
timestamp 1668240031
transform -1 0 31832 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_8  _1840_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1668240031
transform 1 0 27600 0 1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_2  _1841_
timestamp 1668240031
transform -1 0 35144 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1842_
timestamp 1668240031
transform -1 0 34408 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1843_
timestamp 1668240031
transform -1 0 34408 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1844_
timestamp 1668240031
transform -1 0 31464 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1845_
timestamp 1668240031
transform -1 0 28060 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1846_
timestamp 1668240031
transform 1 0 29992 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1847_
timestamp 1668240031
transform 1 0 36340 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1848_
timestamp 1668240031
transform -1 0 31464 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1849_
timestamp 1668240031
transform -1 0 36340 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1850_
timestamp 1668240031
transform 1 0 36340 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1851_
timestamp 1668240031
transform 1 0 27232 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1852_
timestamp 1668240031
transform 1 0 36708 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1853_
timestamp 1668240031
transform -1 0 36616 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1854_
timestamp 1668240031
transform -1 0 35880 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1855_
timestamp 1668240031
transform 1 0 35972 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1856_
timestamp 1668240031
transform -1 0 32568 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1857_
timestamp 1668240031
transform -1 0 31004 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1858_
timestamp 1668240031
transform -1 0 32568 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1859_
timestamp 1668240031
transform -1 0 30636 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1860_
timestamp 1668240031
transform -1 0 29256 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1861_
timestamp 1668240031
transform -1 0 28612 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1862_
timestamp 1668240031
transform 1 0 27232 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1863_
timestamp 1668240031
transform 1 0 29532 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1864_
timestamp 1668240031
transform -1 0 27416 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1865_
timestamp 1668240031
transform -1 0 27416 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1866_
timestamp 1668240031
transform -1 0 27416 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1867_
timestamp 1668240031
transform -1 0 27968 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1868_
timestamp 1668240031
transform -1 0 29624 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1869_
timestamp 1668240031
transform -1 0 28612 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1870_
timestamp 1668240031
transform -1 0 27140 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1871_
timestamp 1668240031
transform 1 0 27508 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1872_
timestamp 1668240031
transform 1 0 27692 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1873_
timestamp 1668240031
transform 1 0 27140 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1874_
timestamp 1668240031
transform 1 0 29164 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1875_
timestamp 1668240031
transform 1 0 27784 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1876_
timestamp 1668240031
transform 1 0 26404 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1877_
timestamp 1668240031
transform -1 0 27324 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1878_
timestamp 1668240031
transform -1 0 26680 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1879_
timestamp 1668240031
transform -1 0 26680 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1880_
timestamp 1668240031
transform -1 0 26588 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1881_
timestamp 1668240031
transform -1 0 27140 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1882_
timestamp 1668240031
transform -1 0 26220 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1883_
timestamp 1668240031
transform -1 0 26864 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1884_
timestamp 1668240031
transform -1 0 22540 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1885_
timestamp 1668240031
transform 1 0 26404 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1886_
timestamp 1668240031
transform 1 0 26404 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1887_
timestamp 1668240031
transform -1 0 20976 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1888_
timestamp 1668240031
transform 1 0 21252 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1889_
timestamp 1668240031
transform 1 0 21804 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1890_
timestamp 1668240031
transform -1 0 17112 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1891_
timestamp 1668240031
transform 1 0 20332 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1892_
timestamp 1668240031
transform 1 0 20056 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1893_
timestamp 1668240031
transform -1 0 16376 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1894_
timestamp 1668240031
transform 1 0 16744 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1895_
timestamp 1668240031
transform -1 0 12420 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1896_
timestamp 1668240031
transform 1 0 13524 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1897_
timestamp 1668240031
transform 1 0 12236 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1898_
timestamp 1668240031
transform 1 0 8372 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1899_
timestamp 1668240031
transform 1 0 7176 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1900_
timestamp 1668240031
transform 1 0 7176 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1901_
timestamp 1668240031
transform 1 0 12880 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1902_
timestamp 1668240031
transform -1 0 13340 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1903_
timestamp 1668240031
transform 1 0 9108 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1904_
timestamp 1668240031
transform 1 0 6532 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1905_
timestamp 1668240031
transform 1 0 6532 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1906_
timestamp 1668240031
transform 1 0 15824 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1907_
timestamp 1668240031
transform -1 0 11960 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1908_
timestamp 1668240031
transform -1 0 11224 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1909_
timestamp 1668240031
transform 1 0 13524 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1910_
timestamp 1668240031
transform 1 0 15180 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1911_
timestamp 1668240031
transform -1 0 20056 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1912_
timestamp 1668240031
transform -1 0 21068 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1913_
timestamp 1668240031
transform -1 0 21344 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1914_
timestamp 1668240031
transform 1 0 21988 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1915_
timestamp 1668240031
transform 1 0 21252 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1916_
timestamp 1668240031
transform 1 0 18676 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1917_
timestamp 1668240031
transform -1 0 17388 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1918_
timestamp 1668240031
transform 1 0 16100 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1919_
timestamp 1668240031
transform 1 0 14260 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1920_
timestamp 1668240031
transform -1 0 15456 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1921_
timestamp 1668240031
transform 1 0 14628 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1922_
timestamp 1668240031
transform -1 0 14536 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1923_
timestamp 1668240031
transform 1 0 12144 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1924_
timestamp 1668240031
transform 1 0 9752 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1925_
timestamp 1668240031
transform 1 0 8372 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1926_
timestamp 1668240031
transform -1 0 7452 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1927_
timestamp 1668240031
transform -1 0 11040 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1928_
timestamp 1668240031
transform -1 0 16376 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1929_
timestamp 1668240031
transform 1 0 11960 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1930_
timestamp 1668240031
transform -1 0 15456 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1931_
timestamp 1668240031
transform 1 0 8096 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1932_
timestamp 1668240031
transform -1 0 7360 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1933_
timestamp 1668240031
transform -1 0 7452 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1934_
timestamp 1668240031
transform -1 0 8004 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1935_
timestamp 1668240031
transform -1 0 6256 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1936_
timestamp 1668240031
transform -1 0 10948 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1937_
timestamp 1668240031
transform 1 0 7728 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1938_
timestamp 1668240031
transform -1 0 10580 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1939_
timestamp 1668240031
transform 1 0 17112 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1940_
timestamp 1668240031
transform -1 0 14444 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1941_
timestamp 1668240031
transform -1 0 14536 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1942_
timestamp 1668240031
transform -1 0 13800 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1943_
timestamp 1668240031
transform 1 0 17204 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1944_
timestamp 1668240031
transform 1 0 16836 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1945_
timestamp 1668240031
transform 1 0 13524 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1946_
timestamp 1668240031
transform -1 0 11224 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1947_
timestamp 1668240031
transform 1 0 11960 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1948_
timestamp 1668240031
transform 1 0 14812 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1949_
timestamp 1668240031
transform 1 0 18584 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1950_
timestamp 1668240031
transform 1 0 28612 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1951_
timestamp 1668240031
transform -1 0 22264 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1952_
timestamp 1668240031
transform -1 0 24840 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1953_
timestamp 1668240031
transform 1 0 30636 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1954_
timestamp 1668240031
transform 1 0 33672 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1955_
timestamp 1668240031
transform -1 0 34960 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1956_
timestamp 1668240031
transform 1 0 33856 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1957_
timestamp 1668240031
transform 1 0 34868 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1958_
timestamp 1668240031
transform 1 0 33764 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1959_
timestamp 1668240031
transform -1 0 31096 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1960_
timestamp 1668240031
transform 1 0 26404 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_8  _1961_
timestamp 1668240031
transform 1 0 29716 0 1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_2  _1962_
timestamp 1668240031
transform -1 0 28612 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1963_
timestamp 1668240031
transform 1 0 28980 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1964_
timestamp 1668240031
transform 1 0 28980 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1965_
timestamp 1668240031
transform 1 0 30360 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1966_
timestamp 1668240031
transform 1 0 29716 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1967_
timestamp 1668240031
transform -1 0 33948 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1968_
timestamp 1668240031
transform 1 0 34868 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1969_
timestamp 1668240031
transform -1 0 33948 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1970_
timestamp 1668240031
transform -1 0 33120 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1971_
timestamp 1668240031
transform -1 0 31832 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1972_
timestamp 1668240031
transform -1 0 32476 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1973_
timestamp 1668240031
transform 1 0 32292 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1974_
timestamp 1668240031
transform -1 0 33856 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1975_
timestamp 1668240031
transform -1 0 33856 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1976_
timestamp 1668240031
transform 1 0 34224 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1977_
timestamp 1668240031
transform -1 0 33212 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1978_
timestamp 1668240031
transform -1 0 33672 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1979_
timestamp 1668240031
transform -1 0 33764 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1980_
timestamp 1668240031
transform -1 0 33304 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1981_
timestamp 1668240031
transform 1 0 32936 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1982_
timestamp 1668240031
transform -1 0 33580 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1983_
timestamp 1668240031
transform -1 0 32568 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1984_
timestamp 1668240031
transform -1 0 32384 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1985_
timestamp 1668240031
transform 1 0 33120 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1986_
timestamp 1668240031
transform -1 0 35144 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1987_
timestamp 1668240031
transform 1 0 35880 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1988_
timestamp 1668240031
transform -1 0 36248 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1989_
timestamp 1668240031
transform 1 0 36616 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1990_
timestamp 1668240031
transform -1 0 33396 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1991_
timestamp 1668240031
transform -1 0 31740 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1992_
timestamp 1668240031
transform -1 0 31832 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1993_
timestamp 1668240031
transform -1 0 33304 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1994_
timestamp 1668240031
transform 1 0 32752 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1995_
timestamp 1668240031
transform -1 0 15640 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1996_
timestamp 1668240031
transform -1 0 14996 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1997_
timestamp 1668240031
transform 1 0 17020 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1998_
timestamp 1668240031
transform -1 0 18032 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1999_
timestamp 1668240031
transform -1 0 17112 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2000_
timestamp 1668240031
transform -1 0 16836 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2001_
timestamp 1668240031
transform 1 0 17204 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2002_
timestamp 1668240031
transform -1 0 16836 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2003_
timestamp 1668240031
transform -1 0 18952 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2004_
timestamp 1668240031
transform -1 0 17756 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _2005_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1668240031
transform 1 0 24656 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2006_
timestamp 1668240031
transform 1 0 24564 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2007_
timestamp 1668240031
transform 1 0 22264 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2008_
timestamp 1668240031
transform 1 0 21988 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2009_
timestamp 1668240031
transform 1 0 21068 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2010_
timestamp 1668240031
transform -1 0 23000 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2011_
timestamp 1668240031
transform 1 0 21620 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2012_
timestamp 1668240031
transform 1 0 21988 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2013_
timestamp 1668240031
transform 1 0 21988 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2014_
timestamp 1668240031
transform 1 0 24564 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2015_
timestamp 1668240031
transform 1 0 22080 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2016_
timestamp 1668240031
transform 1 0 23000 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2017_
timestamp 1668240031
transform 1 0 22724 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2018_
timestamp 1668240031
transform 1 0 22264 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2019_
timestamp 1668240031
transform 1 0 24196 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2020_
timestamp 1668240031
transform 1 0 21988 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2021_
timestamp 1668240031
transform 1 0 22080 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2022_
timestamp 1668240031
transform 1 0 20700 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2023_
timestamp 1668240031
transform 1 0 20424 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2024_
timestamp 1668240031
transform 1 0 20884 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2025_
timestamp 1668240031
transform -1 0 23000 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2026_
timestamp 1668240031
transform 1 0 20700 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2027_
timestamp 1668240031
transform 1 0 21988 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2028_
timestamp 1668240031
transform 1 0 22172 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2029_
timestamp 1668240031
transform 1 0 24196 0 -1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2030_
timestamp 1668240031
transform 1 0 22080 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2031_
timestamp 1668240031
transform 1 0 20608 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2032_
timestamp 1668240031
transform -1 0 19964 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2033_
timestamp 1668240031
transform 1 0 16836 0 -1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2034_
timestamp 1668240031
transform 1 0 16468 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2035_
timestamp 1668240031
transform 1 0 17296 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2036_
timestamp 1668240031
transform 1 0 17112 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2037_
timestamp 1668240031
transform 1 0 13984 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2038_
timestamp 1668240031
transform -1 0 15916 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2039_
timestamp 1668240031
transform 1 0 14260 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2040_
timestamp 1668240031
transform -1 0 14812 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2041_
timestamp 1668240031
transform 1 0 10764 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2042_
timestamp 1668240031
transform 1 0 7820 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2043_
timestamp 1668240031
transform 1 0 7820 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2044_
timestamp 1668240031
transform 1 0 10396 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2045_
timestamp 1668240031
transform 1 0 9752 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2046_
timestamp 1668240031
transform 1 0 9292 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2047_
timestamp 1668240031
transform 1 0 7636 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2048_
timestamp 1668240031
transform 1 0 6532 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2049_
timestamp 1668240031
transform 1 0 7360 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2050_
timestamp 1668240031
transform 1 0 9384 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2051_
timestamp 1668240031
transform 1 0 12328 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2052_
timestamp 1668240031
transform 1 0 14536 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2053_
timestamp 1668240031
transform -1 0 19044 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2054_
timestamp 1668240031
transform -1 0 19780 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2055_
timestamp 1668240031
transform 1 0 17480 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2056_
timestamp 1668240031
transform -1 0 20056 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2057_
timestamp 1668240031
transform -1 0 21528 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2058_
timestamp 1668240031
transform 1 0 19412 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2059_
timestamp 1668240031
transform 1 0 16836 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2060_
timestamp 1668240031
transform 1 0 14536 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2061_
timestamp 1668240031
transform 1 0 12604 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2062_
timestamp 1668240031
transform 1 0 11684 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2063_
timestamp 1668240031
transform 1 0 11684 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2064_
timestamp 1668240031
transform 1 0 10488 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2065_
timestamp 1668240031
transform 1 0 9108 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2066_
timestamp 1668240031
transform 1 0 6624 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2067_
timestamp 1668240031
transform 1 0 6808 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2068_
timestamp 1668240031
transform 1 0 8004 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2069_
timestamp 1668240031
transform 1 0 9384 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2070_
timestamp 1668240031
transform 1 0 11224 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2071_
timestamp 1668240031
transform 1 0 9108 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2072_
timestamp 1668240031
transform 1 0 6532 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2073_
timestamp 1668240031
transform 1 0 6256 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2074_
timestamp 1668240031
transform 1 0 6532 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2075_
timestamp 1668240031
transform -1 0 9292 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2076_
timestamp 1668240031
transform -1 0 11224 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2077_
timestamp 1668240031
transform 1 0 8464 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2078_
timestamp 1668240031
transform 1 0 8280 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2079_
timestamp 1668240031
transform 1 0 10304 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2080_
timestamp 1668240031
transform 1 0 10120 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2081_
timestamp 1668240031
transform 1 0 11684 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2082_
timestamp 1668240031
transform 1 0 14260 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2083_
timestamp 1668240031
transform -1 0 15364 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2084_
timestamp 1668240031
transform 1 0 11776 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2085_
timestamp 1668240031
transform 1 0 11316 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2086_
timestamp 1668240031
transform 1 0 10488 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2087_
timestamp 1668240031
transform -1 0 16376 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2088_
timestamp 1668240031
transform 1 0 17112 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2089_
timestamp 1668240031
transform 1 0 19320 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2090_
timestamp 1668240031
transform 1 0 21988 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2091_
timestamp 1668240031
transform 1 0 27232 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2092_
timestamp 1668240031
transform 1 0 30912 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2093_
timestamp 1668240031
transform 1 0 31004 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2094_
timestamp 1668240031
transform 1 0 29992 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2095_
timestamp 1668240031
transform 1 0 32016 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2096_
timestamp 1668240031
transform 1 0 31924 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2097_
timestamp 1668240031
transform -1 0 31648 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2098_
timestamp 1668240031
transform 1 0 28704 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2099_
timestamp 1668240031
transform 1 0 26220 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2100_
timestamp 1668240031
transform -1 0 30820 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _2101_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1668240031
transform 1 0 35236 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2102_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1668240031
transform -1 0 32016 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2103_
timestamp 1668240031
transform 1 0 34868 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2104_
timestamp 1668240031
transform -1 0 36524 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2105_
timestamp 1668240031
transform -1 0 36984 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2106_
timestamp 1668240031
transform 1 0 35052 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2107_
timestamp 1668240031
transform -1 0 34408 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2108_
timestamp 1668240031
transform 1 0 34960 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2109_
timestamp 1668240031
transform 1 0 30176 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2110_
timestamp 1668240031
transform -1 0 31648 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2111_
timestamp 1668240031
transform -1 0 29900 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2112_
timestamp 1668240031
transform -1 0 28980 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2113_
timestamp 1668240031
transform -1 0 28888 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2114_
timestamp 1668240031
transform 1 0 24932 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2115_
timestamp 1668240031
transform 1 0 24840 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2116_
timestamp 1668240031
transform 1 0 24932 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2117_
timestamp 1668240031
transform -1 0 27416 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2118_
timestamp 1668240031
transform 1 0 25484 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2119_
timestamp 1668240031
transform 1 0 26404 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2120_
timestamp 1668240031
transform 1 0 27140 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2121_
timestamp 1668240031
transform 1 0 26680 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2122_
timestamp 1668240031
transform 1 0 27140 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2123_
timestamp 1668240031
transform 1 0 27140 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2124_
timestamp 1668240031
transform 1 0 27140 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2125_
timestamp 1668240031
transform 1 0 26588 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2126_
timestamp 1668240031
transform 1 0 27140 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2127_
timestamp 1668240031
transform 1 0 27140 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2128_
timestamp 1668240031
transform 1 0 24932 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2129_
timestamp 1668240031
transform 1 0 24840 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2130_
timestamp 1668240031
transform 1 0 24932 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2131_
timestamp 1668240031
transform 1 0 24656 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2132_
timestamp 1668240031
transform 1 0 24656 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2133_
timestamp 1668240031
transform 1 0 24840 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2134_
timestamp 1668240031
transform 1 0 24932 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2135_
timestamp 1668240031
transform 1 0 24932 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2136_
timestamp 1668240031
transform 1 0 24840 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2137_
timestamp 1668240031
transform 1 0 19412 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2138_
timestamp 1668240031
transform 1 0 20240 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2139_
timestamp 1668240031
transform 1 0 21988 0 -1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2140_
timestamp 1668240031
transform 1 0 15732 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2141_
timestamp 1668240031
transform 1 0 19412 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2142_
timestamp 1668240031
transform 1 0 19044 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2143_
timestamp 1668240031
transform -1 0 17756 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2144_
timestamp 1668240031
transform 1 0 15824 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2145_
timestamp 1668240031
transform 1 0 13800 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2146_
timestamp 1668240031
transform 1 0 11684 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2147_
timestamp 1668240031
transform 1 0 9108 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2148_
timestamp 1668240031
transform 1 0 6624 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2149_
timestamp 1668240031
transform 1 0 6716 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2150_
timestamp 1668240031
transform 1 0 12236 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2151_
timestamp 1668240031
transform 1 0 11960 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2152_
timestamp 1668240031
transform 1 0 11132 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2153_
timestamp 1668240031
transform 1 0 6440 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2154_
timestamp 1668240031
transform 1 0 6532 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _2155_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1668240031
transform 1 0 10212 0 1 27200
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _2156_
timestamp 1668240031
transform 1 0 11776 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2157_
timestamp 1668240031
transform 1 0 13248 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2158_
timestamp 1668240031
transform 1 0 15824 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2159_
timestamp 1668240031
transform 1 0 18676 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2160_
timestamp 1668240031
transform 1 0 19688 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2161_
timestamp 1668240031
transform 1 0 19688 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2162_
timestamp 1668240031
transform 1 0 20332 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2163_
timestamp 1668240031
transform 1 0 20424 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2164_
timestamp 1668240031
transform -1 0 21252 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2165_
timestamp 1668240031
transform 1 0 16836 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2166_
timestamp 1668240031
transform 1 0 14536 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2167_
timestamp 1668240031
transform 1 0 14076 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2168_
timestamp 1668240031
transform 1 0 14260 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2169_
timestamp 1668240031
transform 1 0 12972 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2170_
timestamp 1668240031
transform 1 0 11132 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2171_
timestamp 1668240031
transform 1 0 9200 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2172_
timestamp 1668240031
transform 1 0 7452 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2173_
timestamp 1668240031
transform 1 0 6992 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2174_
timestamp 1668240031
transform 1 0 9384 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2175_
timestamp 1668240031
transform 1 0 11316 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2176_
timestamp 1668240031
transform 1 0 13248 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2177_
timestamp 1668240031
transform 1 0 9108 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2178_
timestamp 1668240031
transform 1 0 5980 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2179_
timestamp 1668240031
transform 1 0 6072 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2180_
timestamp 1668240031
transform 1 0 6072 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2181_
timestamp 1668240031
transform -1 0 8372 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2182_
timestamp 1668240031
transform 1 0 9108 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2183_
timestamp 1668240031
transform 1 0 6808 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2184_
timestamp 1668240031
transform 1 0 8924 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2185_
timestamp 1668240031
transform 1 0 12052 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2186_
timestamp 1668240031
transform 1 0 11776 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2187_
timestamp 1668240031
transform 1 0 12144 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2188_
timestamp 1668240031
transform 1 0 16836 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2189_
timestamp 1668240031
transform 1 0 15824 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2190_
timestamp 1668240031
transform -1 0 15640 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2191_
timestamp 1668240031
transform -1 0 13524 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2192_
timestamp 1668240031
transform 1 0 12328 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2193_
timestamp 1668240031
transform -1 0 16376 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2194_
timestamp 1668240031
transform 1 0 17112 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2195_
timestamp 1668240031
transform 1 0 20240 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2196_
timestamp 1668240031
transform -1 0 25116 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2197_
timestamp 1668240031
transform 1 0 29716 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2198_
timestamp 1668240031
transform 1 0 32660 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2199_
timestamp 1668240031
transform 1 0 32752 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2200_
timestamp 1668240031
transform 1 0 32844 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2201_
timestamp 1668240031
transform 1 0 33028 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2202_
timestamp 1668240031
transform 1 0 32752 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2203_
timestamp 1668240031
transform 1 0 29716 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2204_
timestamp 1668240031
transform 1 0 26864 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2205_
timestamp 1668240031
transform 1 0 26036 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2206_
timestamp 1668240031
transform -1 0 30820 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _2207_
timestamp 1668240031
transform -1 0 31832 0 1 23936
box -38 -48 2154 592
use sky130_fd_sc_hd__dfstp_1  _2208_
timestamp 1668240031
transform 1 0 29716 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_1  _2209_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1668240031
transform -1 0 34500 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2210_
timestamp 1668240031
transform 1 0 33396 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2211_
timestamp 1668240031
transform -1 0 32568 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _2212_
timestamp 1668240031
transform 1 0 30912 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2213_
timestamp 1668240031
transform 1 0 31280 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2214_
timestamp 1668240031
transform -1 0 32844 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2215_
timestamp 1668240031
transform -1 0 32660 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2216_
timestamp 1668240031
transform 1 0 31280 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2217_
timestamp 1668240031
transform 1 0 32292 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2218_
timestamp 1668240031
transform -1 0 33028 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2219_
timestamp 1668240031
transform -1 0 34132 0 -1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2220_
timestamp 1668240031
transform -1 0 31832 0 -1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2221_
timestamp 1668240031
transform 1 0 31004 0 1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2222_
timestamp 1668240031
transform 1 0 32292 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2223_
timestamp 1668240031
transform 1 0 33764 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2224_
timestamp 1668240031
transform 1 0 34868 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2225_
timestamp 1668240031
transform 1 0 33856 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2226_
timestamp 1668240031
transform 1 0 35328 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2227_
timestamp 1668240031
transform -1 0 34408 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2228_
timestamp 1668240031
transform 1 0 30360 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2229_
timestamp 1668240031
transform 1 0 29992 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2230_
timestamp 1668240031
transform 1 0 29992 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2231_
timestamp 1668240031
transform -1 0 34132 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2232_
timestamp 1668240031
transform 1 0 14260 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2233_
timestamp 1668240031
transform 1 0 13892 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2234_
timestamp 1668240031
transform -1 0 18676 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2235_
timestamp 1668240031
transform 1 0 16560 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2236_
timestamp 1668240031
transform -1 0 17480 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2237_
timestamp 1668240031
transform -1 0 16192 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2238_
timestamp 1668240031
transform -1 0 18676 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2239_
timestamp 1668240031
transform -1 0 17756 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2240_
timestamp 1668240031
transform -1 0 19964 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2241_
timestamp 1668240031
transform 1 0 16284 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk_in pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1668240031
transform -1 0 21436 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_ref_in
timestamp 1668240031
transform -1 0 35328 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_vco_in
timestamp 1668240031
transform 1 0 32292 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_ref_in
timestamp 1668240031
transform -1 0 33028 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_vco_in
timestamp 1668240031
transform -1 0 30452 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_ref_in
timestamp 1668240031
transform -1 0 33028 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_vco_in
timestamp 1668240031
transform 1 0 32292 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_clk_in
timestamp 1668240031
transform 1 0 12788 0 1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_clk_in
timestamp 1668240031
transform -1 0 16284 0 1 6528
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_clk_in
timestamp 1668240031
transform -1 0 12696 0 -1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_clk_in
timestamp 1668240031
transform 1 0 12696 0 1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_clk_in
timestamp 1668240031
transform 1 0 25024 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_clk_in
timestamp 1668240031
transform 1 0 27508 0 1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_clk_in
timestamp 1668240031
transform 1 0 23184 0 -1 15232
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_clk_in
timestamp 1668240031
transform 1 0 25668 0 -1 15232
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_clk_in
timestamp 1668240031
transform -1 0 10948 0 1 23936
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_clk_in
timestamp 1668240031
transform 1 0 11960 0 1 23936
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_clk_in
timestamp 1668240031
transform -1 0 10856 0 1 30464
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_clk_in
timestamp 1668240031
transform 1 0 12328 0 -1 31552
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_clk_in
timestamp 1668240031
transform 1 0 20240 0 -1 27200
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_clk_in
timestamp 1668240031
transform 1 0 22816 0 -1 27200
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_clk_in
timestamp 1668240031
transform -1 0 20516 0 -1 33728
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_clk_in
timestamp 1668240031
transform 1 0 21804 0 1 32640
box -38 -48 1050 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input1 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1668240031
transform 1 0 32292 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  input2
timestamp 1668240031
transform 1 0 29716 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1668240031
transform 1 0 25208 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1668240031
transform 1 0 34868 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output5
timestamp 1668240031
transform -1 0 36984 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output6
timestamp 1668240031
transform -1 0 37168 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output7
timestamp 1668240031
transform -1 0 37168 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output8
timestamp 1668240031
transform 1 0 1748 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output9
timestamp 1668240031
transform 1 0 4692 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output10
timestamp 1668240031
transform 1 0 7636 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output11
timestamp 1668240031
transform -1 0 9936 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output12
timestamp 1668240031
transform -1 0 11224 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output13
timestamp 1668240031
transform -1 0 16376 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output14
timestamp 1668240031
transform -1 0 19320 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output15
timestamp 1668240031
transform 1 0 22356 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output16
timestamp 1668240031
transform -1 0 36984 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output17
timestamp 1668240031
transform 1 0 1564 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output18
timestamp 1668240031
transform 1 0 1564 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output19
timestamp 1668240031
transform 1 0 1564 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output20
timestamp 1668240031
transform 1 0 1564 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output21
timestamp 1668240031
transform 1 0 1564 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output22
timestamp 1668240031
transform 1 0 1564 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output23
timestamp 1668240031
transform 1 0 1564 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output24
timestamp 1668240031
transform 1 0 1564 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output25
timestamp 1668240031
transform 1 0 1564 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output26
timestamp 1668240031
transform 1 0 1564 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output27
timestamp 1668240031
transform 1 0 1564 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output28
timestamp 1668240031
transform 1 0 21252 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output29
timestamp 1668240031
transform 1 0 19412 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output30
timestamp 1668240031
transform -1 0 11960 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output31
timestamp 1668240031
transform -1 0 10580 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output32
timestamp 1668240031
transform 1 0 9660 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output33
timestamp 1668240031
transform 1 0 6992 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output34
timestamp 1668240031
transform 1 0 4232 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output35
timestamp 1668240031
transform 1 0 1564 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output36
timestamp 1668240031
transform -1 0 36984 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output37
timestamp 1668240031
transform -1 0 37168 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output38
timestamp 1668240031
transform -1 0 36984 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output39
timestamp 1668240031
transform -1 0 37168 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output40
timestamp 1668240031
transform -1 0 37168 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output41
timestamp 1668240031
transform -1 0 36984 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output42
timestamp 1668240031
transform -1 0 37168 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output43
timestamp 1668240031
transform -1 0 37168 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  wrapper_44 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1668240031
transform -1 0 26128 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  wrapper_45
timestamp 1668240031
transform -1 0 30820 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  wrapper_46
timestamp 1668240031
transform -1 0 34408 0 1 38080
box -38 -48 314 592
<< labels >>
flabel metal2 s 26238 0 26294 800 0 FreeSans 224 90 0 0 clk_in
port 0 nsew signal input
flabel metal3 s 37949 38632 38749 38752 0 FreeSans 480 0 0 0 corner[0]
port 1 nsew signal tristate
flabel metal3 s 37949 34960 38749 35080 0 FreeSans 480 0 0 0 corner[1]
port 2 nsew signal tristate
flabel metal3 s 37949 31288 38749 31408 0 FreeSans 480 0 0 0 corner[2]
port 3 nsew signal tristate
flabel metal2 s 1674 40093 1730 40893 0 FreeSans 224 90 0 0 dac[0]
port 4 nsew signal tristate
flabel metal2 s 4618 40093 4674 40893 0 FreeSans 224 90 0 0 dac[1]
port 5 nsew signal tristate
flabel metal2 s 7562 40093 7618 40893 0 FreeSans 224 90 0 0 dac[2]
port 6 nsew signal tristate
flabel metal2 s 10506 40093 10562 40893 0 FreeSans 224 90 0 0 dac[3]
port 7 nsew signal tristate
flabel metal2 s 13450 40093 13506 40893 0 FreeSans 224 90 0 0 dac[4]
port 8 nsew signal tristate
flabel metal2 s 16394 40093 16450 40893 0 FreeSans 224 90 0 0 dac[5]
port 9 nsew signal tristate
flabel metal2 s 19338 40093 19394 40893 0 FreeSans 224 90 0 0 dac[6]
port 10 nsew signal tristate
flabel metal2 s 22282 40093 22338 40893 0 FreeSans 224 90 0 0 dac[7]
port 11 nsew signal tristate
flabel metal2 s 25226 40093 25282 40893 0 FreeSans 224 90 0 0 dac[8]
port 12 nsew signal tristate
flabel metal2 s 28170 40093 28226 40893 0 FreeSans 224 90 0 0 dac[9]
port 13 nsew signal tristate
flabel metal2 s 31758 0 31814 800 0 FreeSans 224 90 0 0 load
port 14 nsew signal input
flabel metal2 s 34058 40093 34114 40893 0 FreeSans 224 90 0 0 lock
port 15 nsew signal tristate
flabel metal2 s 28998 0 29054 800 0 FreeSans 224 90 0 0 read
port 16 nsew signal input
flabel metal2 s 37002 40093 37058 40893 0 FreeSans 224 90 0 0 ref_in
port 17 nsew signal input
flabel metal2 s 23478 0 23534 800 0 FreeSans 224 90 0 0 reset
port 18 nsew signal input
flabel metal2 s 34518 0 34574 800 0 FreeSans 224 90 0 0 s_in
port 19 nsew signal input
flabel metal2 s 37278 0 37334 800 0 FreeSans 224 90 0 0 s_out
port 20 nsew signal tristate
flabel metal3 s 0 34960 800 35080 0 FreeSans 480 0 0 0 slope_ctrl[0]
port 21 nsew signal tristate
flabel metal3 s 0 38632 800 38752 0 FreeSans 480 0 0 0 slope_ctrl[1]
port 22 nsew signal tristate
flabel metal3 s 0 31288 800 31408 0 FreeSans 480 0 0 0 slope_ctrl[2]
port 23 nsew signal tristate
flabel metal3 s 0 1912 800 2032 0 FreeSans 480 0 0 0 vbias1[0]
port 24 nsew signal tristate
flabel metal3 s 0 5584 800 5704 0 FreeSans 480 0 0 0 vbias1[1]
port 25 nsew signal tristate
flabel metal3 s 0 9256 800 9376 0 FreeSans 480 0 0 0 vbias1[2]
port 26 nsew signal tristate
flabel metal3 s 0 12928 800 13048 0 FreeSans 480 0 0 0 vbias1[3]
port 27 nsew signal tristate
flabel metal3 s 0 16600 800 16720 0 FreeSans 480 0 0 0 vbias1[4]
port 28 nsew signal tristate
flabel metal3 s 0 20272 800 20392 0 FreeSans 480 0 0 0 vbias1[5]
port 29 nsew signal tristate
flabel metal3 s 0 23944 800 24064 0 FreeSans 480 0 0 0 vbias1[6]
port 30 nsew signal tristate
flabel metal3 s 0 27616 800 27736 0 FreeSans 480 0 0 0 vbias1[7]
port 31 nsew signal tristate
flabel metal2 s 20718 0 20774 800 0 FreeSans 224 90 0 0 vbias2[0]
port 32 nsew signal tristate
flabel metal2 s 17958 0 18014 800 0 FreeSans 224 90 0 0 vbias2[1]
port 33 nsew signal tristate
flabel metal2 s 15198 0 15254 800 0 FreeSans 224 90 0 0 vbias2[2]
port 34 nsew signal tristate
flabel metal2 s 12438 0 12494 800 0 FreeSans 224 90 0 0 vbias2[3]
port 35 nsew signal tristate
flabel metal2 s 9678 0 9734 800 0 FreeSans 224 90 0 0 vbias2[4]
port 36 nsew signal tristate
flabel metal2 s 6918 0 6974 800 0 FreeSans 224 90 0 0 vbias2[5]
port 37 nsew signal tristate
flabel metal2 s 4158 0 4214 800 0 FreeSans 224 90 0 0 vbias2[6]
port 38 nsew signal tristate
flabel metal2 s 1398 0 1454 800 0 FreeSans 224 90 0 0 vbias2[7]
port 39 nsew signal tristate
flabel metal3 s 37949 1912 38749 2032 0 FreeSans 480 0 0 0 vbias3[0]
port 40 nsew signal tristate
flabel metal3 s 37949 5584 38749 5704 0 FreeSans 480 0 0 0 vbias3[1]
port 41 nsew signal tristate
flabel metal3 s 37949 9256 38749 9376 0 FreeSans 480 0 0 0 vbias3[2]
port 42 nsew signal tristate
flabel metal3 s 37949 12928 38749 13048 0 FreeSans 480 0 0 0 vbias3[3]
port 43 nsew signal tristate
flabel metal3 s 37949 16600 38749 16720 0 FreeSans 480 0 0 0 vbias3[4]
port 44 nsew signal tristate
flabel metal3 s 37949 20272 38749 20392 0 FreeSans 480 0 0 0 vbias3[5]
port 45 nsew signal tristate
flabel metal3 s 37949 23944 38749 24064 0 FreeSans 480 0 0 0 vbias3[6]
port 46 nsew signal tristate
flabel metal3 s 37949 27616 38749 27736 0 FreeSans 480 0 0 0 vbias3[7]
port 47 nsew signal tristate
flabel metal2 s 31114 40093 31170 40893 0 FreeSans 224 90 0 0 vco_in
port 48 nsew signal input
flabel metal4 s 4208 2128 4528 38672 0 FreeSans 1920 90 0 0 vdd
port 49 nsew power bidirectional
flabel metal4 s 34928 2128 35248 38672 0 FreeSans 1920 90 0 0 vdd
port 49 nsew power bidirectional
flabel metal5 s 1056 5346 37676 5666 0 FreeSans 2560 0 0 0 vdd
port 49 nsew power bidirectional
flabel metal5 s 1056 35982 37676 36302 0 FreeSans 2560 0 0 0 vdd
port 49 nsew power bidirectional
flabel metal4 s 4868 2128 5188 38672 0 FreeSans 1920 90 0 0 vss
port 50 nsew ground bidirectional
flabel metal4 s 35588 2128 35908 38672 0 FreeSans 1920 90 0 0 vss
port 50 nsew ground bidirectional
flabel metal5 s 1056 6006 37676 6326 0 FreeSans 2560 0 0 0 vss
port 50 nsew ground bidirectional
flabel metal5 s 1056 36642 37676 36962 0 FreeSans 2560 0 0 0 vss
port 50 nsew ground bidirectional
rlabel metal1 19366 38624 19366 38624 0 vdd
rlabel metal1 19366 38080 19366 38080 0 vss
rlabel metal1 30544 24582 30544 24582 0 _0000_
rlabel metal1 31832 30770 31832 30770 0 _0001_
rlabel metal1 31326 30158 31326 30158 0 _0002_
rlabel metal2 33074 32674 33074 32674 0 _0003_
rlabel metal2 32430 33762 32430 33762 0 _0004_
rlabel metal2 30314 35258 30314 35258 0 _0005_
rlabel metal1 32108 35734 32108 35734 0 _0006_
rlabel metal2 32706 34850 32706 34850 0 _0007_
rlabel metal2 33810 37604 33810 37604 0 _0008_
rlabel metal2 31510 38046 31510 38046 0 _0009_
rlabel metal1 30314 36686 30314 36686 0 _0010_
rlabel metal1 32982 17102 32982 17102 0 _0011_
rlabel metal1 34040 17850 34040 17850 0 _0012_
rlabel metal1 35236 17238 35236 17238 0 _0013_
rlabel metal2 34270 14756 34270 14756 0 _0014_
rlabel metal1 35512 14586 35512 14586 0 _0015_
rlabel metal1 33258 14586 33258 14586 0 _0016_
rlabel metal2 30682 15708 30682 15708 0 _0017_
rlabel metal2 30314 17374 30314 17374 0 _0018_
rlabel metal2 30314 18462 30314 18462 0 _0019_
rlabel metal2 31050 19108 31050 19108 0 _0020_
rlabel metal2 26082 9146 26082 9146 0 _0021_
rlabel metal2 25530 9792 25530 9792 0 _0022_
rlabel metal1 23736 9622 23736 9622 0 _0023_
rlabel metal2 23046 11560 23046 11560 0 _0024_
rlabel metal1 22310 12614 22310 12614 0 _0025_
rlabel metal1 21482 14042 21482 14042 0 _0026_
rlabel metal2 22678 15266 22678 15266 0 _0027_
rlabel metal2 22770 17374 22770 17374 0 _0028_
rlabel metal2 22954 18462 22954 18462 0 _0029_
rlabel metal1 24840 18394 24840 18394 0 _0030_
rlabel metal2 24334 20366 24334 20366 0 _0031_
rlabel metal2 24702 21182 24702 21182 0 _0032_
rlabel metal2 23690 22168 23690 22168 0 _0033_
rlabel metal1 23460 22066 23460 22066 0 _0034_
rlabel metal2 25898 24990 25898 24990 0 _0035_
rlabel metal2 23690 24582 23690 24582 0 _0036_
rlabel metal2 25346 26112 25346 26112 0 _0037_
rlabel metal2 22126 27098 22126 27098 0 _0038_
rlabel metal2 23506 28016 23506 28016 0 _0039_
rlabel metal1 21528 29274 21528 29274 0 _0040_
rlabel metal2 21390 30872 21390 30872 0 _0041_
rlabel metal1 21436 32198 21436 32198 0 _0042_
rlabel metal1 22533 33558 22533 33558 0 _0043_
rlabel metal1 25714 34680 25714 34680 0 _0044_
rlabel metal1 24833 37910 24833 37910 0 _0045_
rlabel metal2 23138 37502 23138 37502 0 _0046_
rlabel metal2 22034 35258 22034 35258 0 _0047_
rlabel metal2 19182 36312 19182 36312 0 _0048_
rlabel metal1 17940 36278 17940 36278 0 _0049_
rlabel metal1 18407 34986 18407 34986 0 _0050_
rlabel metal1 17979 33558 17979 33558 0 _0051_
rlabel metal1 18354 32198 18354 32198 0 _0052_
rlabel metal2 15272 32334 15272 32334 0 _0053_
rlabel metal2 11086 32606 11086 32606 0 _0054_
rlabel metal2 15594 34850 15594 34850 0 _0055_
rlabel metal2 12374 34782 12374 34782 0 _0056_
rlabel metal2 12098 36312 12098 36312 0 _0057_
rlabel metal2 9154 36142 9154 36142 0 _0058_
rlabel metal1 8142 32470 8142 32470 0 _0059_
rlabel metal1 11132 34510 11132 34510 0 _0060_
rlabel metal1 10488 32198 10488 32198 0 _0061_
rlabel metal1 10021 29206 10021 29206 0 _0062_
rlabel metal2 9246 31790 9246 31790 0 _0063_
rlabel metal2 7314 27846 7314 27846 0 _0064_
rlabel metal1 8464 26554 8464 26554 0 _0065_
rlabel metal1 9515 28118 9515 28118 0 _0066_
rlabel metal2 13662 29342 13662 29342 0 _0067_
rlabel metal2 15594 28968 15594 28968 0 _0068_
rlabel metal1 18913 29206 18913 29206 0 _0069_
rlabel metal1 19189 27030 19189 27030 0 _0070_
rlabel metal1 18584 23290 18584 23290 0 _0071_
rlabel metal2 19274 21998 19274 21998 0 _0072_
rlabel metal1 20424 16218 20424 16218 0 _0073_
rlabel metal1 19964 16218 19964 16218 0 _0074_
rlabel metal1 18124 16218 18124 16218 0 _0075_
rlabel metal1 15640 16218 15640 16218 0 _0076_
rlabel metal1 13195 18326 13195 18326 0 _0077_
rlabel metal2 12466 20264 12466 20264 0 _0078_
rlabel metal1 12236 22066 12236 22066 0 _0079_
rlabel metal2 12098 22338 12098 22338 0 _0080_
rlabel metal2 10074 22372 10074 22372 0 _0081_
rlabel metal2 8050 22338 8050 22338 0 _0082_
rlabel metal1 7912 21318 7912 21318 0 _0083_
rlabel metal1 9292 19686 9292 19686 0 _0084_
rlabel metal1 9890 17850 9890 17850 0 _0085_
rlabel metal1 11868 16422 11868 16422 0 _0086_
rlabel metal1 10212 16218 10212 16218 0 _0087_
rlabel metal1 6617 17238 6617 17238 0 _0088_
rlabel metal1 6325 15334 6325 15334 0 _0089_
rlabel metal2 7130 13022 7130 13022 0 _0090_
rlabel metal1 8563 7446 8563 7446 0 _0091_
rlabel metal1 10580 8058 10580 8058 0 _0092_
rlabel metal2 9522 10846 9522 10846 0 _0093_
rlabel metal1 8786 13430 8786 13430 0 _0094_
rlabel metal1 12128 13226 12128 13226 0 _0095_
rlabel metal1 10764 12070 10764 12070 0 _0096_
rlabel metal2 12098 9112 12098 9112 0 _0097_
rlabel metal1 14168 8806 14168 8806 0 _0098_
rlabel metal2 14398 7582 14398 7582 0 _0099_
rlabel metal1 12880 7174 12880 7174 0 _0100_
rlabel metal1 11868 5338 11868 5338 0 _0101_
rlabel metal1 10672 4998 10672 4998 0 _0102_
rlabel metal2 15502 4590 15502 4590 0 _0103_
rlabel metal1 18262 4998 18262 4998 0 _0104_
rlabel metal1 20608 4454 20608 4454 0 _0105_
rlabel metal1 23598 3706 23598 3706 0 _0106_
rlabel metal2 28106 3944 28106 3944 0 _0107_
rlabel metal1 32660 4794 32660 4794 0 _0108_
rlabel metal1 33212 6834 33212 6834 0 _0109_
rlabel metal2 31694 9112 31694 9112 0 _0110_
rlabel metal1 34277 11050 34277 11050 0 _0111_
rlabel metal1 33863 13226 33863 13226 0 _0112_
rlabel metal1 33994 10778 33994 10778 0 _0113_
rlabel metal1 30820 7514 30820 7514 0 _0114_
rlabel metal1 27837 6698 27837 6698 0 _0115_
rlabel metal1 30084 5882 30084 5882 0 _0116_
rlabel metal2 36478 25534 36478 25534 0 _0117_
rlabel metal1 31280 24786 31280 24786 0 _0118_
rlabel metal2 36202 27846 36202 27846 0 _0119_
rlabel metal1 36386 25466 36386 25466 0 _0120_
rlabel metal1 35413 23018 35413 23018 0 _0121_
rlabel metal2 36478 23222 36478 23222 0 _0122_
rlabel metal1 34691 19754 34691 19754 0 _0123_
rlabel metal1 36064 21862 36064 21862 0 _0124_
rlabel metal2 31602 20740 31602 20740 0 _0125_
rlabel metal2 30866 19618 30866 19618 0 _0126_
rlabel metal1 29263 10710 29263 10710 0 _0127_
rlabel metal1 28389 12138 28389 12138 0 _0128_
rlabel metal1 28159 13226 28159 13226 0 _0129_
rlabel metal1 27922 11866 27922 11866 0 _0130_
rlabel metal1 28021 13974 28021 13974 0 _0131_
rlabel metal2 27278 13634 27278 13634 0 _0132_
rlabel metal2 26634 15640 26634 15640 0 _0133_
rlabel metal1 27055 16490 27055 16490 0 _0134_
rlabel metal2 27830 17102 27830 17102 0 _0135_
rlabel metal1 29079 19414 29079 19414 0 _0136_
rlabel metal1 28251 19754 28251 19754 0 _0137_
rlabel metal1 27455 21590 27455 21590 0 _0138_
rlabel metal1 27784 22066 27784 22066 0 _0139_
rlabel metal1 27876 23290 27876 23290 0 _0140_
rlabel metal1 28711 25194 28711 25194 0 _0141_
rlabel metal2 27922 25364 27922 25364 0 _0142_
rlabel metal1 27048 27846 27048 27846 0 _0143_
rlabel metal1 27048 26554 27048 26554 0 _0144_
rlabel metal2 26542 28968 26542 28968 0 _0145_
rlabel metal1 26503 29546 26503 29546 0 _0146_
rlabel metal1 26319 31382 26319 31382 0 _0147_
rlabel metal1 26549 31790 26549 31790 0 _0148_
rlabel metal1 26174 33082 26174 33082 0 _0149_
rlabel metal1 26680 33082 26680 33082 0 _0150_
rlabel metal1 26503 37162 26503 37162 0 _0151_
rlabel metal2 26542 35870 26542 35870 0 _0152_
rlabel metal2 20838 34374 20838 34374 0 _0153_
rlabel metal1 21344 36890 21344 36890 0 _0154_
rlabel metal2 22770 37128 22770 37128 0 _0155_
rlabel metal1 17020 36346 17020 36346 0 _0156_
rlabel metal2 20470 32674 20470 32674 0 _0157_
rlabel metal1 20286 31790 20286 31790 0 _0158_
rlabel metal1 16330 30294 16330 30294 0 _0159_
rlabel metal2 16882 33320 16882 33320 0 _0160_
rlabel metal2 15226 37502 15226 37502 0 _0161_
rlabel metal2 12374 37638 12374 37638 0 _0162_
rlabel metal1 8878 37094 8878 37094 0 _0163_
rlabel metal1 7360 36006 7360 36006 0 _0164_
rlabel metal2 7314 32402 7314 32402 0 _0165_
rlabel metal2 13018 34238 13018 34238 0 _0166_
rlabel metal2 13386 32266 13386 32266 0 _0167_
rlabel metal1 9890 29546 9890 29546 0 _0168_
rlabel metal2 6578 31110 6578 31110 0 _0169_
rlabel metal2 7314 29342 7314 29342 0 _0170_
rlabel metal1 11783 27370 11783 27370 0 _0171_
rlabel metal1 11270 26758 11270 26758 0 _0172_
rlabel metal1 13839 27030 13839 27030 0 _0173_
rlabel metal1 15955 27370 15955 27370 0 _0174_
rlabel metal1 19964 28390 19964 28390 0 _0175_
rlabel metal1 20976 25466 20976 25466 0 _0176_
rlabel metal1 21160 24038 21160 24038 0 _0177_
rlabel metal1 21949 21998 21949 21998 0 _0178_
rlabel metal1 21344 20230 21344 20230 0 _0179_
rlabel metal2 18814 19176 18814 19176 0 _0180_
rlabel metal1 17158 16422 17158 16422 0 _0181_
rlabel metal1 14858 18938 14858 18938 0 _0182_
rlabel metal1 15364 20774 15364 20774 0 _0183_
rlabel metal1 14904 21658 14904 21658 0 _0184_
rlabel metal2 14398 23868 14398 23868 0 _0185_
rlabel metal1 12236 25670 12236 25670 0 _0186_
rlabel metal1 9936 24786 9936 24786 0 _0187_
rlabel metal2 8510 25262 8510 25262 0 _0188_
rlabel metal1 7537 23766 7537 23766 0 _0189_
rlabel metal1 10856 20774 10856 20774 0 _0190_
rlabel metal2 12098 17816 12098 17816 0 _0191_
rlabel metal1 15226 15130 15226 15130 0 _0192_
rlabel metal1 9062 18394 9062 18394 0 _0193_
rlabel metal1 7268 18394 7268 18394 0 _0194_
rlabel metal1 7360 13498 7360 13498 0 _0195_
rlabel metal1 7643 9962 7643 9962 0 _0196_
rlabel metal1 6479 8534 6479 8534 0 _0197_
rlabel metal2 10810 9554 10810 9554 0 _0198_
rlabel metal2 7866 12002 7866 12002 0 _0199_
rlabel metal1 10396 15334 10396 15334 0 _0200_
rlabel metal1 14030 12954 14030 12954 0 _0201_
rlabel metal1 13853 12138 13853 12138 0 _0202_
rlabel metal1 13616 11050 13616 11050 0 _0203_
rlabel metal1 17756 8058 17756 8058 0 _0204_
rlabel metal1 16928 6086 16928 6086 0 _0205_
rlabel metal2 13662 4998 13662 4998 0 _0206_
rlabel metal1 11539 2346 11539 2346 0 _0207_
rlabel metal2 13110 3298 13110 3298 0 _0208_
rlabel metal2 14950 2822 14950 2822 0 _0209_
rlabel metal2 18722 2856 18722 2856 0 _0210_
rlabel metal1 22034 2618 22034 2618 0 _0211_
rlabel metal1 24525 3094 24525 3094 0 _0212_
rlabel metal2 30774 4318 30774 4318 0 _0213_
rlabel metal1 33764 5338 33764 5338 0 _0214_
rlabel metal2 34822 7888 34822 7888 0 _0215_
rlabel metal1 33948 9146 33948 9146 0 _0216_
rlabel metal2 35006 11934 35006 11934 0 _0217_
rlabel metal2 33810 13294 33810 13294 0 _0218_
rlabel metal2 31050 13736 31050 13736 0 _0219_
rlabel metal1 27094 8602 27094 8602 0 _0220_
rlabel metal1 27975 5678 27975 5678 0 _0221_
rlabel metal2 29118 6120 29118 6120 0 _0222_
rlabel metal1 29755 24174 29755 24174 0 _0223_
rlabel metal2 30498 23528 30498 23528 0 _0224_
rlabel metal1 33081 30634 33081 30634 0 _0225_
rlabel metal1 33219 31790 33219 31790 0 _0226_
rlabel metal1 33212 32470 33212 32470 0 _0227_
rlabel metal2 33074 33728 33074 33728 0 _0228_
rlabel metal1 33304 35258 33304 35258 0 _0229_
rlabel metal1 33672 36006 33672 36006 0 _0230_
rlabel metal2 33166 34544 33166 34544 0 _0231_
rlabel metal2 33074 38046 33074 38046 0 _0232_
rlabel metal2 33442 37604 33442 37604 0 _0233_
rlabel metal2 32430 37706 32430 37706 0 _0234_
rlabel metal2 33258 16898 33258 16898 0 _0235_
rlabel metal1 35052 18598 35052 18598 0 _0236_
rlabel metal1 35972 16762 35972 16762 0 _0237_
rlabel metal2 36110 15470 36110 15470 0 _0238_
rlabel metal2 36754 15674 36754 15674 0 _0239_
rlabel metal1 33166 15130 33166 15130 0 _0240_
rlabel metal2 31786 15028 31786 15028 0 _0241_
rlabel metal2 31694 16898 31694 16898 0 _0242_
rlabel metal1 32246 18292 32246 18292 0 _0243_
rlabel metal1 32844 18938 32844 18938 0 _0244_
rlabel metal1 15410 24786 15410 24786 0 _0245_
rlabel metal1 15042 24718 15042 24718 0 _0246_
rlabel metal1 17204 26758 17204 26758 0 _0247_
rlabel metal1 17940 24650 17940 24650 0 _0248_
rlabel metal1 16836 23834 16836 23834 0 _0249_
rlabel metal1 15555 23018 15555 23018 0 _0250_
rlabel metal2 17342 22814 17342 22814 0 _0251_
rlabel metal2 16698 21352 16698 21352 0 _0252_
rlabel metal1 18860 18938 18860 18938 0 _0253_
rlabel metal2 17618 19992 17618 19992 0 _0254_
rlabel metal1 25162 8058 25162 8058 0 _0255_
rlabel metal1 24840 9418 24840 9418 0 _0256_
rlabel metal2 22586 10200 22586 10200 0 _0257_
rlabel metal2 22310 11492 22310 11492 0 _0258_
rlabel metal1 21436 12138 21436 12138 0 _0259_
rlabel metal1 22678 14280 22678 14280 0 _0260_
rlabel metal2 21942 15708 21942 15708 0 _0261_
rlabel metal2 22310 16932 22310 16932 0 _0262_
rlabel metal1 22448 17850 22448 17850 0 _0263_
rlabel metal1 24472 18666 24472 18666 0 _0264_
rlabel metal2 22402 19822 22402 19822 0 _0265_
rlabel metal2 24610 20196 24610 20196 0 _0266_
rlabel metal1 23460 21862 23460 21862 0 _0267_
rlabel metal2 22586 23528 22586 23528 0 _0268_
rlabel metal1 25024 24718 25024 24718 0 _0269_
rlabel metal2 22310 24990 22310 24990 0 _0270_
rlabel metal1 23506 25806 23506 25806 0 _0271_
rlabel metal2 21022 26520 21022 26520 0 _0272_
rlabel metal1 20884 28186 20884 28186 0 _0273_
rlabel metal2 21206 29784 21206 29784 0 _0274_
rlabel metal1 23046 30634 23046 30634 0 _0275_
rlabel metal1 21521 31994 21521 31994 0 _0276_
rlabel metal1 22494 32538 22494 32538 0 _0277_
rlabel metal1 22632 34646 22632 34646 0 _0278_
rlabel metal2 24518 38046 24518 38046 0 _0279_
rlabel metal2 22402 36958 22402 36958 0 _0280_
rlabel metal2 20930 35224 20930 35224 0 _0281_
rlabel metal1 19642 36856 19642 36856 0 _0282_
rlabel metal2 17158 38046 17158 38046 0 _0283_
rlabel metal2 16330 34850 16330 34850 0 _0284_
rlabel metal2 17618 33694 17618 33694 0 _0285_
rlabel metal1 17250 31450 17250 31450 0 _0286_
rlabel metal1 12167 31450 12167 31450 0 _0287_
rlabel metal1 15048 32198 15048 32198 0 _0288_
rlabel metal1 14168 34986 14168 34986 0 _0289_
rlabel metal1 15327 34374 15327 34374 0 _0290_
rlabel metal1 11040 36074 11040 36074 0 _0291_
rlabel metal1 7774 35598 7774 35598 0 _0292_
rlabel metal1 7774 32538 7774 32538 0 _0293_
rlabel metal2 10718 34204 10718 34204 0 _0294_
rlabel metal1 9384 31858 9384 31858 0 _0295_
rlabel metal1 8878 29206 8878 29206 0 _0296_
rlabel metal1 7590 31382 7590 31382 0 _0297_
rlabel metal2 6854 28254 6854 28254 0 _0298_
rlabel metal2 7774 26724 7774 26724 0 _0299_
rlabel metal1 10718 27982 10718 27982 0 _0300_
rlabel metal2 12650 28900 12650 28900 0 _0301_
rlabel metal1 15088 29070 15088 29070 0 _0302_
rlabel metal1 19053 28934 19053 28934 0 _0303_
rlabel metal1 20056 27030 20056 27030 0 _0304_
rlabel metal2 17802 23902 17802 23902 0 _0305_
rlabel metal1 19688 20026 19688 20026 0 _0306_
rlabel metal2 21206 17374 21206 17374 0 _0307_
rlabel metal1 19228 16218 19228 16218 0 _0308_
rlabel metal2 17158 16354 17158 16354 0 _0309_
rlabel metal1 15042 15674 15042 15674 0 _0310_
rlabel metal2 12926 18734 12926 18734 0 _0311_
rlabel metal1 11822 20502 11822 20502 0 _0312_
rlabel metal1 11960 22678 11960 22678 0 _0313_
rlabel metal2 10810 22610 10810 22610 0 _0314_
rlabel metal1 9476 22202 9476 22202 0 _0315_
rlabel metal1 7130 22202 7130 22202 0 _0316_
rlabel metal1 7268 20570 7268 20570 0 _0317_
rlabel metal1 8372 19278 8372 19278 0 _0318_
rlabel metal1 9338 18190 9338 18190 0 _0319_
rlabel metal1 11352 15674 11352 15674 0 _0320_
rlabel metal1 8786 16218 8786 16218 0 _0321_
rlabel metal2 6854 17153 6854 17153 0 _0322_
rlabel metal1 6302 15130 6302 15130 0 _0323_
rlabel metal1 6624 12410 6624 12410 0 _0324_
rlabel metal2 8970 7582 8970 7582 0 _0325_
rlabel metal2 10902 8670 10902 8670 0 _0326_
rlabel metal2 8786 11118 8786 11118 0 _0327_
rlabel metal2 8602 14110 8602 14110 0 _0328_
rlabel metal2 10626 13532 10626 13532 0 _0329_
rlabel metal1 10580 10778 10580 10778 0 _0330_
rlabel metal1 11592 9486 11592 9486 0 _0331_
rlabel metal1 14122 8602 14122 8602 0 _0332_
rlabel metal1 15042 7480 15042 7480 0 _0333_
rlabel metal1 12137 6970 12137 6970 0 _0334_
rlabel metal2 11638 5916 11638 5916 0 _0335_
rlabel metal2 10810 3944 10810 3944 0 _0336_
rlabel metal1 15778 2618 15778 2618 0 _0337_
rlabel metal2 17526 3876 17526 3876 0 _0338_
rlabel metal2 19642 4318 19642 4318 0 _0339_
rlabel metal1 22172 4182 22172 4182 0 _0340_
rlabel metal2 27554 4318 27554 4318 0 _0341_
rlabel metal1 31602 4794 31602 4794 0 _0342_
rlabel metal1 33113 8058 33113 8058 0 _0343_
rlabel metal1 30360 9622 30360 9622 0 _0344_
rlabel metal1 32844 10234 32844 10234 0 _0345_
rlabel metal2 31694 13464 31694 13464 0 _0346_
rlabel metal1 32669 11322 32669 11322 0 _0347_
rlabel metal1 29992 8398 29992 8398 0 _0348_
rlabel metal1 26857 6970 26857 6970 0 _0349_
rlabel metal1 30866 6426 30866 6426 0 _0350_
rlabel metal2 35650 26588 35650 26588 0 _0351_
rlabel metal2 31694 26588 31694 26588 0 _0352_
rlabel metal2 35190 28254 35190 28254 0 _0353_
rlabel metal1 36064 25466 36064 25466 0 _0354_
rlabel metal1 35972 22746 35972 22746 0 _0355_
rlabel metal1 35006 23630 35006 23630 0 _0356_
rlabel metal2 34086 20060 34086 20060 0 _0357_
rlabel metal1 35282 20570 35282 20570 0 _0358_
rlabel metal1 30590 20570 30590 20570 0 _0359_
rlabel metal2 31326 19992 31326 19992 0 _0360_
rlabel metal2 29578 11390 29578 11390 0 _0361_
rlabel metal1 28796 10234 28796 10234 0 _0362_
rlabel metal2 28842 13090 28842 13090 0 _0363_
rlabel metal2 24058 11730 24058 11730 0 _0364_
rlabel metal1 24978 13974 24978 13974 0 _0365_
rlabel metal1 24656 13430 24656 13430 0 _0366_
rlabel metal1 27738 15130 27738 15130 0 _0367_
rlabel metal1 25290 16762 25290 16762 0 _0368_
rlabel metal2 26726 17884 26726 17884 0 _0369_
rlabel metal2 27002 19108 27002 19108 0 _0370_
rlabel metal2 27002 20060 27002 20060 0 _0371_
rlabel metal1 27048 21454 27048 21454 0 _0372_
rlabel metal1 27462 22712 27462 22712 0 _0373_
rlabel metal1 27002 23290 27002 23290 0 _0374_
rlabel metal1 27048 24922 27048 24922 0 _0375_
rlabel metal1 27600 25942 27600 25942 0 _0376_
rlabel metal1 26956 27098 26956 27098 0 _0377_
rlabel metal1 25438 27098 25438 27098 0 _0378_
rlabel metal1 25484 28730 25484 28730 0 _0379_
rlabel metal2 25254 30124 25254 30124 0 _0380_
rlabel metal1 24610 31382 24610 31382 0 _0381_
rlabel metal2 24978 32028 24978 32028 0 _0382_
rlabel metal1 24794 33422 24794 33422 0 _0383_
rlabel metal1 25760 34034 25760 34034 0 _0384_
rlabel metal2 25254 37740 25254 37740 0 _0385_
rlabel metal2 25162 35870 25162 35870 0 _0386_
rlabel metal2 18262 34272 18262 34272 0 _0387_
rlabel metal1 20562 37128 20562 37128 0 _0388_
rlabel metal1 22310 37944 22310 37944 0 _0389_
rlabel metal1 16100 36890 16100 36890 0 _0390_
rlabel metal1 19320 32810 19320 32810 0 _0391_
rlabel metal2 19458 30974 19458 30974 0 _0392_
rlabel metal1 17112 32198 17112 32198 0 _0393_
rlabel metal1 15630 33082 15630 33082 0 _0394_
rlabel metal2 14122 37502 14122 37502 0 _0395_
rlabel metal1 11592 36890 11592 36890 0 _0396_
rlabel metal2 9430 37468 9430 37468 0 _0397_
rlabel metal2 6762 35360 6762 35360 0 _0398_
rlabel metal2 7038 33116 7038 33116 0 _0399_
rlabel metal1 12190 33558 12190 33558 0 _0400_
rlabel metal1 11720 31994 11720 31994 0 _0401_
rlabel metal1 11270 29682 11270 29682 0 _0402_
rlabel metal1 6716 30634 6716 30634 0 _0403_
rlabel metal1 6486 29206 6486 29206 0 _0404_
rlabel metal1 10166 27370 10166 27370 0 _0405_
rlabel metal1 12006 26418 12006 26418 0 _0406_
rlabel metal2 13570 27710 13570 27710 0 _0407_
rlabel via1 16139 27642 16139 27642 0 _0408_
rlabel metal1 18998 28152 18998 28152 0 _0409_
rlabel metal1 19642 25942 19642 25942 0 _0410_
rlabel metal2 20010 24174 20010 24174 0 _0411_
rlabel metal1 19918 21896 19918 21896 0 _0412_
rlabel metal2 20746 19992 20746 19992 0 _0413_
rlabel metal1 16652 18122 16652 18122 0 _0414_
rlabel metal1 15686 16456 15686 16456 0 _0415_
rlabel metal2 13754 19108 13754 19108 0 _0416_
rlabel metal1 14444 20502 14444 20502 0 _0417_
rlabel metal1 14342 22202 14342 22202 0 _0418_
rlabel metal2 13294 23902 13294 23902 0 _0419_
rlabel metal1 11454 25160 11454 25160 0 _0420_
rlabel metal2 8602 25636 8602 25636 0 _0421_
rlabel metal2 7774 24990 7774 24990 0 _0422_
rlabel metal2 7314 23460 7314 23460 0 _0423_
rlabel metal1 9844 20502 9844 20502 0 _0424_
rlabel metal1 11684 17578 11684 17578 0 _0425_
rlabel metal2 13570 16286 13570 16286 0 _0426_
rlabel metal1 8326 17850 8326 17850 0 _0427_
rlabel metal2 6026 18530 6026 18530 0 _0428_
rlabel metal1 6026 14314 6026 14314 0 _0429_
rlabel metal2 6394 10472 6394 10472 0 _0430_
rlabel metal1 6026 8364 6026 8364 0 _0431_
rlabel metal1 9016 9962 9016 9962 0 _0432_
rlabel metal1 7406 11322 7406 11322 0 _0433_
rlabel metal1 8878 14926 8878 14926 0 _0434_
rlabel metal1 12144 13974 12144 13974 0 _0435_
rlabel metal1 12098 12104 12098 12104 0 _0436_
rlabel metal2 11822 10404 11822 10404 0 _0437_
rlabel metal2 17158 8228 17158 8228 0 _0438_
rlabel metal2 16146 6188 16146 6188 0 _0439_
rlabel metal2 15318 5440 15318 5440 0 _0440_
rlabel metal1 13064 2346 13064 2346 0 _0441_
rlabel metal1 12650 3128 12650 3128 0 _0442_
rlabel metal2 16882 4046 16882 4046 0 _0443_
rlabel metal2 17434 2788 17434 2788 0 _0444_
rlabel metal2 19918 3298 19918 3298 0 _0445_
rlabel metal2 24794 2788 24794 2788 0 _0446_
rlabel metal1 29532 4658 29532 4658 0 _0447_
rlabel metal1 33948 6222 33948 6222 0 _0448_
rlabel metal1 33534 6630 33534 6630 0 _0449_
rlabel metal1 33304 9622 33304 9622 0 _0450_
rlabel metal1 32936 10778 32936 10778 0 _0451_
rlabel metal2 33074 13566 33074 13566 0 _0452_
rlabel metal1 30038 13192 30038 13192 0 _0453_
rlabel metal2 27186 8466 27186 8466 0 _0454_
rlabel metal2 26358 5916 26358 5916 0 _0455_
rlabel metal1 31050 5338 31050 5338 0 _0456_
rlabel metal1 34561 29206 34561 29206 0 _0457_
rlabel metal2 33074 30022 33074 30022 0 _0458_
rlabel metal1 32353 28458 32353 28458 0 _0459_
rlabel metal1 29486 15674 29486 15674 0 _0460_
rlabel metal1 30222 16422 30222 16422 0 _0461_
rlabel metal1 30222 29172 30222 29172 0 _0462_
rlabel metal1 29348 34510 29348 34510 0 _0463_
rlabel metal1 29210 33830 29210 33830 0 _0464_
rlabel metal1 28106 29716 28106 29716 0 _0465_
rlabel metal2 27922 29852 27922 29852 0 _0466_
rlabel metal1 27646 30736 27646 30736 0 _0467_
rlabel metal1 27324 30362 27324 30362 0 _0468_
rlabel metal1 27784 29614 27784 29614 0 _0469_
rlabel metal1 28704 29818 28704 29818 0 _0470_
rlabel metal2 28382 29580 28382 29580 0 _0471_
rlabel metal1 29164 29274 29164 29274 0 _0472_
rlabel metal1 29624 37230 29624 37230 0 _0473_
rlabel metal1 29532 27846 29532 27846 0 _0474_
rlabel metal1 28612 27982 28612 27982 0 _0475_
rlabel metal1 29716 28730 29716 28730 0 _0476_
rlabel metal1 28704 28594 28704 28594 0 _0477_
rlabel metal1 28520 28186 28520 28186 0 _0478_
rlabel metal2 29026 29206 29026 29206 0 _0479_
rlabel metal1 29440 29546 29440 29546 0 _0480_
rlabel metal2 29578 29444 29578 29444 0 _0481_
rlabel metal1 29716 25874 29716 25874 0 _0482_
rlabel metal2 30406 25466 30406 25466 0 _0483_
rlabel metal2 31786 25636 31786 25636 0 _0484_
rlabel metal1 31050 25738 31050 25738 0 _0485_
rlabel metal1 28980 24922 28980 24922 0 _0486_
rlabel metal1 29072 23290 29072 23290 0 _0487_
rlabel metal1 29900 24650 29900 24650 0 _0488_
rlabel metal1 29854 25908 29854 25908 0 _0489_
rlabel metal1 29578 25262 29578 25262 0 _0490_
rlabel metal1 35052 24242 35052 24242 0 _0491_
rlabel metal1 31510 20468 31510 20468 0 _0492_
rlabel metal2 30314 21862 30314 21862 0 _0493_
rlabel metal2 30866 20876 30866 20876 0 _0494_
rlabel metal1 32706 20876 32706 20876 0 _0495_
rlabel metal1 33304 20910 33304 20910 0 _0496_
rlabel metal2 33718 21284 33718 21284 0 _0497_
rlabel metal1 34684 20910 34684 20910 0 _0498_
rlabel metal2 35006 20604 35006 20604 0 _0499_
rlabel metal1 33856 20366 33856 20366 0 _0500_
rlabel metal1 34362 20434 34362 20434 0 _0501_
rlabel metal1 34684 25194 34684 25194 0 _0502_
rlabel metal2 33626 23834 33626 23834 0 _0503_
rlabel metal1 34224 23630 34224 23630 0 _0504_
rlabel metal2 34454 23868 34454 23868 0 _0505_
rlabel metal1 35098 25296 35098 25296 0 _0506_
rlabel metal2 34822 25024 34822 25024 0 _0507_
rlabel metal1 35512 22610 35512 22610 0 _0508_
rlabel metal1 34224 25874 34224 25874 0 _0509_
rlabel metal1 33718 26010 33718 26010 0 _0510_
rlabel metal2 34270 26758 34270 26758 0 _0511_
rlabel metal2 35512 25874 35512 25874 0 _0512_
rlabel metal1 34592 27438 34592 27438 0 _0513_
rlabel metal1 35558 27642 35558 27642 0 _0514_
rlabel metal1 34592 28186 34592 28186 0 _0515_
rlabel metal1 32338 27540 32338 27540 0 _0516_
rlabel metal2 30774 27200 30774 27200 0 _0517_
rlabel metal1 31372 26962 31372 26962 0 _0518_
rlabel metal1 24794 11220 24794 11220 0 _0519_
rlabel metal2 30958 5066 30958 5066 0 _0520_
rlabel metal1 30268 5338 30268 5338 0 _0521_
rlabel metal1 30682 6630 30682 6630 0 _0522_
rlabel metal2 28474 6528 28474 6528 0 _0523_
rlabel metal1 27278 6426 27278 6426 0 _0524_
rlabel metal1 29486 7854 29486 7854 0 _0525_
rlabel metal1 30820 8058 30820 8058 0 _0526_
rlabel metal1 30222 10778 30222 10778 0 _0527_
rlabel metal1 31372 11594 31372 11594 0 _0528_
rlabel metal1 31510 12410 31510 12410 0 _0529_
rlabel metal1 21850 2958 21850 2958 0 _0530_
rlabel metal2 31510 13430 31510 13430 0 _0531_
rlabel metal1 32108 11866 32108 11866 0 _0532_
rlabel metal1 32660 10030 32660 10030 0 _0533_
rlabel metal1 31970 8942 31970 8942 0 _0534_
rlabel metal2 31418 9894 31418 9894 0 _0535_
rlabel metal1 33120 8602 33120 8602 0 _0536_
rlabel metal1 34868 7854 34868 7854 0 _0537_
rlabel metal2 32890 5984 32890 5984 0 _0538_
rlabel metal2 32154 4794 32154 4794 0 _0539_
rlabel metal1 28888 4590 28888 4590 0 _0540_
rlabel metal1 27968 4590 27968 4590 0 _0541_
rlabel metal1 24794 4080 24794 4080 0 _0542_
rlabel metal1 23782 3978 23782 3978 0 _0543_
rlabel metal1 22172 4590 22172 4590 0 _0544_
rlabel metal1 21482 3094 21482 3094 0 _0545_
rlabel metal1 20194 3162 20194 3162 0 _0546_
rlabel metal1 18308 3706 18308 3706 0 _0547_
rlabel metal1 17894 3502 17894 3502 0 _0548_
rlabel metal1 16284 3706 16284 3706 0 _0549_
rlabel metal1 15824 2414 15824 2414 0 _0550_
rlabel metal1 13156 3978 13156 3978 0 _0551_
rlabel metal1 13892 6222 13892 6222 0 _0552_
rlabel metal1 10672 4590 10672 4590 0 _0553_
rlabel metal1 12742 4250 12742 4250 0 _0554_
rlabel metal1 12098 4794 12098 4794 0 _0555_
rlabel metal1 13202 5338 13202 5338 0 _0556_
rlabel metal1 12512 6426 12512 6426 0 _0557_
rlabel metal2 14674 5882 14674 5882 0 _0558_
rlabel metal1 15502 5882 15502 5882 0 _0559_
rlabel metal1 14812 8058 14812 8058 0 _0560_
rlabel metal1 13800 8466 13800 8466 0 _0561_
rlabel metal1 12834 8942 12834 8942 0 _0562_
rlabel metal1 11546 9146 11546 9146 0 _0563_
rlabel metal1 8050 9010 8050 9010 0 _0564_
rlabel metal2 12374 11526 12374 11526 0 _0565_
rlabel metal1 11040 10642 11040 10642 0 _0566_
rlabel metal2 10810 13600 10810 13600 0 _0567_
rlabel metal1 10488 12954 10488 12954 0 _0568_
rlabel metal1 9430 13294 9430 13294 0 _0569_
rlabel metal1 8786 13498 8786 13498 0 _0570_
rlabel metal1 9292 11866 9292 11866 0 _0571_
rlabel metal1 8740 11730 8740 11730 0 _0572_
rlabel metal2 9890 9146 9890 9146 0 _0573_
rlabel metal2 9660 16796 9660 16796 0 _0574_
rlabel metal1 11546 8976 11546 8976 0 _0575_
rlabel metal1 7452 8874 7452 8874 0 _0576_
rlabel metal1 7682 7854 7682 7854 0 _0577_
rlabel metal1 6992 9418 6992 9418 0 _0578_
rlabel metal1 6394 11866 6394 11866 0 _0579_
rlabel metal2 7038 14518 7038 14518 0 _0580_
rlabel metal1 6256 14994 6256 14994 0 _0581_
rlabel metal1 6762 17578 6762 17578 0 _0582_
rlabel metal1 6164 17646 6164 17646 0 _0583_
rlabel metal1 9476 16150 9476 16150 0 _0584_
rlabel metal1 8280 16082 8280 16082 0 _0585_
rlabel metal1 12006 23596 12006 23596 0 _0586_
rlabel metal2 12282 16320 12282 16320 0 _0587_
rlabel metal1 11362 16082 11362 16082 0 _0588_
rlabel metal1 11132 17306 11132 17306 0 _0589_
rlabel metal1 9706 17510 9706 17510 0 _0590_
rlabel metal2 10626 19584 10626 19584 0 _0591_
rlabel metal1 9430 19482 9430 19482 0 _0592_
rlabel metal1 8556 20570 8556 20570 0 _0593_
rlabel metal1 7820 20434 7820 20434 0 _0594_
rlabel metal1 7314 23018 7314 23018 0 _0595_
rlabel metal2 9798 23426 9798 23426 0 _0596_
rlabel metal2 7498 22474 7498 22474 0 _0597_
rlabel metal1 9476 23834 9476 23834 0 _0598_
rlabel metal2 9338 22746 9338 22746 0 _0599_
rlabel metal2 10810 24208 10810 24208 0 _0600_
rlabel metal2 10626 22746 10626 22746 0 _0601_
rlabel metal1 12834 23086 12834 23086 0 _0602_
rlabel metal2 11362 23732 11362 23732 0 _0603_
rlabel metal1 12512 21862 12512 21862 0 _0604_
rlabel metal1 11776 20910 11776 20910 0 _0605_
rlabel metal1 13570 19482 13570 19482 0 _0606_
rlabel metal1 12374 19414 12374 19414 0 _0607_
rlabel metal1 15916 18802 15916 18802 0 _0608_
rlabel metal1 15042 17646 15042 17646 0 _0609_
rlabel metal2 15410 16490 15410 16490 0 _0610_
rlabel metal1 17434 17306 17434 17306 0 _0611_
rlabel metal2 16974 16524 16974 16524 0 _0612_
rlabel metal2 18906 17408 18906 17408 0 _0613_
rlabel metal2 18906 16524 18906 16524 0 _0614_
rlabel metal2 20378 17850 20378 17850 0 _0615_
rlabel metal1 21068 17646 21068 17646 0 _0616_
rlabel metal1 19596 21658 19596 21658 0 _0617_
rlabel metal1 11178 28526 11178 28526 0 _0618_
rlabel metal2 18906 20842 18906 20842 0 _0619_
rlabel metal1 19320 23290 19320 23290 0 _0620_
rlabel metal2 18354 24378 18354 24378 0 _0621_
rlabel metal1 18998 25466 18998 25466 0 _0622_
rlabel metal2 18906 26962 18906 26962 0 _0623_
rlabel metal1 18722 27574 18722 27574 0 _0624_
rlabel metal2 20286 29308 20286 29308 0 _0625_
rlabel metal1 16514 28730 16514 28730 0 _0626_
rlabel metal2 15778 30022 15778 30022 0 _0627_
rlabel metal1 15042 28186 15042 28186 0 _0628_
rlabel metal1 10350 28594 10350 28594 0 _0629_
rlabel metal1 9798 35156 9798 35156 0 _0630_
rlabel metal1 11868 28186 11868 28186 0 _0631_
rlabel metal2 11914 28220 11914 28220 0 _0632_
rlabel metal1 10718 27098 10718 27098 0 _0633_
rlabel metal2 7958 26826 7958 26826 0 _0634_
rlabel metal1 8648 28458 8648 28458 0 _0635_
rlabel metal1 7498 28526 7498 28526 0 _0636_
rlabel metal1 7636 30090 7636 30090 0 _0637_
rlabel metal2 7038 30702 7038 30702 0 _0638_
rlabel metal2 10166 29818 10166 29818 0 _0639_
rlabel metal1 13018 35564 13018 35564 0 _0640_
rlabel metal1 7866 29614 7866 29614 0 _0641_
rlabel metal1 11270 31450 11270 31450 0 _0642_
rlabel metal1 9706 31450 9706 31450 0 _0643_
rlabel metal1 12236 33082 12236 33082 0 _0644_
rlabel metal1 10350 34612 10350 34612 0 _0645_
rlabel metal1 9568 33082 9568 33082 0 _0646_
rlabel metal1 7590 32402 7590 32402 0 _0647_
rlabel metal2 8878 34816 8878 34816 0 _0648_
rlabel metal1 7866 34714 7866 34714 0 _0649_
rlabel metal1 11270 35530 11270 35530 0 _0650_
rlabel metal1 10994 35802 10994 35802 0 _0651_
rlabel metal1 19964 36210 19964 36210 0 _0652_
rlabel metal1 13156 35802 13156 35802 0 _0653_
rlabel metal1 16330 35700 16330 35700 0 _0654_
rlabel metal1 15456 35802 15456 35802 0 _0655_
rlabel metal2 13570 35292 13570 35292 0 _0656_
rlabel metal1 15042 32912 15042 32912 0 _0657_
rlabel metal1 14490 33082 14490 33082 0 _0658_
rlabel metal2 15594 31178 15594 31178 0 _0659_
rlabel metal2 11914 31110 11914 31110 0 _0660_
rlabel metal1 18308 31450 18308 31450 0 _0661_
rlabel metal1 18538 37298 18538 37298 0 _0662_
rlabel metal1 17204 31314 17204 31314 0 _0663_
rlabel metal1 18860 32538 18860 32538 0 _0664_
rlabel metal1 17802 33082 17802 33082 0 _0665_
rlabel metal1 17986 34714 17986 34714 0 _0666_
rlabel metal2 16422 35020 16422 35020 0 _0667_
rlabel metal2 18170 37264 18170 37264 0 _0668_
rlabel metal1 17572 38318 17572 38318 0 _0669_
rlabel metal1 18998 37230 18998 37230 0 _0670_
rlabel metal1 20562 36788 20562 36788 0 _0671_
rlabel metal1 20332 35802 20332 35802 0 _0672_
rlabel metal1 20884 35666 20884 35666 0 _0673_
rlabel metal1 23874 32946 23874 32946 0 _0674_
rlabel metal1 23460 35802 23460 35802 0 _0675_
rlabel metal2 23046 36788 23046 36788 0 _0676_
rlabel metal1 24012 36890 24012 36890 0 _0677_
rlabel metal1 24426 37434 24426 37434 0 _0678_
rlabel metal1 24748 34986 24748 34986 0 _0679_
rlabel metal2 23322 35462 23322 35462 0 _0680_
rlabel metal1 23828 33966 23828 33966 0 _0681_
rlabel metal2 22862 33116 22862 33116 0 _0682_
rlabel metal1 23276 31790 23276 31790 0 _0683_
rlabel metal1 23046 31858 23046 31858 0 _0684_
rlabel metal1 22586 31994 22586 31994 0 _0685_
rlabel metal1 23092 31450 23092 31450 0 _0686_
rlabel metal2 23598 30906 23598 30906 0 _0687_
rlabel metal2 23506 29818 23506 29818 0 _0688_
rlabel metal1 22770 29818 22770 29818 0 _0689_
rlabel metal1 23184 29274 23184 29274 0 _0690_
rlabel metal2 22126 28492 22126 28492 0 _0691_
rlabel metal1 22908 27438 22908 27438 0 _0692_
rlabel metal2 22218 27132 22218 27132 0 _0693_
rlabel metal1 23736 26350 23736 26350 0 _0694_
rlabel metal1 24380 26350 24380 26350 0 _0695_
rlabel metal1 25714 21454 25714 21454 0 _0696_
rlabel metal1 24104 25262 24104 25262 0 _0697_
rlabel metal1 23000 25262 23000 25262 0 _0698_
rlabel metal2 24978 25466 24978 25466 0 _0699_
rlabel metal1 26220 24786 26220 24786 0 _0700_
rlabel metal2 24426 23936 24426 23936 0 _0701_
rlabel metal1 23598 23834 23598 23834 0 _0702_
rlabel metal2 25346 22848 25346 22848 0 _0703_
rlabel metal1 24518 22066 24518 22066 0 _0704_
rlabel metal2 24978 21114 24978 21114 0 _0705_
rlabel metal1 25990 11730 25990 11730 0 _0706_
rlabel metal2 24794 20298 24794 20298 0 _0707_
rlabel metal1 24058 19822 24058 19822 0 _0708_
rlabel metal1 22954 20026 22954 20026 0 _0709_
rlabel metal1 25392 19482 25392 19482 0 _0710_
rlabel metal1 23920 18734 23920 18734 0 _0711_
rlabel metal1 24242 17578 24242 17578 0 _0712_
rlabel metal1 23000 17646 23000 17646 0 _0713_
rlabel metal1 23828 16558 23828 16558 0 _0714_
rlabel metal1 22586 16558 22586 16558 0 _0715_
rlabel metal1 23828 16218 23828 16218 0 _0716_
rlabel metal1 22724 16082 22724 16082 0 _0717_
rlabel metal1 22908 14042 22908 14042 0 _0718_
rlabel metal1 22862 13804 22862 13804 0 _0719_
rlabel metal1 23046 12954 23046 12954 0 _0720_
rlabel metal1 22011 13294 22011 13294 0 _0721_
rlabel metal1 24058 12206 24058 12206 0 _0722_
rlabel metal1 22494 11152 22494 11152 0 _0723_
rlabel metal2 25346 11526 25346 11526 0 _0724_
rlabel metal1 22770 10676 22770 10676 0 _0725_
rlabel metal2 26266 10880 26266 10880 0 _0726_
rlabel metal2 24978 9996 24978 9996 0 _0727_
rlabel metal1 28382 9486 28382 9486 0 _0728_
rlabel metal2 26358 8602 26358 8602 0 _0729_
rlabel metal1 34454 33082 34454 33082 0 _0730_
rlabel metal2 34362 31110 34362 31110 0 _0731_
rlabel metal1 33350 31314 33350 31314 0 _0732_
rlabel metal1 13570 25874 13570 25874 0 _0733_
rlabel metal1 15042 27098 15042 27098 0 _0734_
rlabel metal1 16468 26350 16468 26350 0 _0735_
rlabel metal1 16146 25840 16146 25840 0 _0736_
rlabel metal1 16698 24786 16698 24786 0 _0737_
rlabel metal1 20976 22950 20976 22950 0 _0738_
rlabel metal1 21988 21386 21988 21386 0 _0739_
rlabel metal1 16882 20468 16882 20468 0 _0740_
rlabel metal1 18952 20434 18952 20434 0 _0741_
rlabel metal1 16284 19482 16284 19482 0 _0742_
rlabel metal1 13524 37978 13524 37978 0 _0743_
rlabel metal1 6095 37842 6095 37842 0 _0744_
rlabel metal1 9062 36890 9062 36890 0 _0745_
rlabel metal2 10350 36550 10350 36550 0 _0746_
rlabel metal2 10488 37094 10488 37094 0 _0747_
rlabel metal1 15456 37842 15456 37842 0 _0748_
rlabel metal1 15088 38318 15088 38318 0 _0749_
rlabel metal1 11730 37842 11730 37842 0 _0750_
rlabel metal1 33166 32300 33166 32300 0 _0751_
rlabel metal1 32982 32368 32982 32368 0 _0752_
rlabel metal1 32522 33422 32522 33422 0 _0753_
rlabel metal1 32039 33490 32039 33490 0 _0754_
rlabel metal1 30866 35598 30866 35598 0 _0755_
rlabel via1 30954 34714 30954 34714 0 _0756_
rlabel metal1 31280 35462 31280 35462 0 _0757_
rlabel metal2 31694 35292 31694 35292 0 _0758_
rlabel metal2 30130 37434 30130 37434 0 _0759_
rlabel metal1 30225 36890 30225 36890 0 _0760_
rlabel metal1 35328 16762 35328 16762 0 _0761_
rlabel metal1 35420 17646 35420 17646 0 _0762_
rlabel metal1 34086 14416 34086 14416 0 _0763_
rlabel metal1 34454 14382 34454 14382 0 _0764_
rlabel metal1 35742 14382 35742 14382 0 _0765_
rlabel metal1 32246 14416 32246 14416 0 _0766_
rlabel metal2 32430 15130 32430 15130 0 _0767_
rlabel metal1 32614 18224 32614 18224 0 _0768_
rlabel metal1 30866 16116 30866 16116 0 _0769_
rlabel metal2 30774 17782 30774 17782 0 _0770_
rlabel metal2 31326 18394 31326 18394 0 _0771_
rlabel metal2 22586 3366 22586 3366 0 _0772_
rlabel metal1 20148 20774 20148 20774 0 _0773_
rlabel metal1 22908 11118 22908 11118 0 _0774_
rlabel metal2 23598 21250 23598 21250 0 _0775_
rlabel metal2 21390 33881 21390 33881 0 _0776_
rlabel metal1 17756 34578 17756 34578 0 _0777_
rlabel metal2 8786 28934 8786 28934 0 _0778_
rlabel metal2 12190 20672 12190 20672 0 _0779_
rlabel metal2 17894 11186 17894 11186 0 _0780_
rlabel metal1 5980 17170 5980 17170 0 _0781_
rlabel metal1 10074 12206 10074 12206 0 _0782_
rlabel metal1 23920 3502 23920 3502 0 _0783_
rlabel metal2 36386 25024 36386 25024 0 _0784_
rlabel metal1 30590 12240 30590 12240 0 _0785_
rlabel metal1 27278 16082 27278 16082 0 _0786_
rlabel metal1 26588 32402 26588 32402 0 _0787_
rlabel metal1 21850 36108 21850 36108 0 _0788_
rlabel metal1 12282 38284 12282 38284 0 _0789_
rlabel metal1 11822 29138 11822 29138 0 _0790_
rlabel metal1 10994 20944 10994 20944 0 _0791_
rlabel metal1 8142 18292 8142 18292 0 _0792_
rlabel metal1 17158 2448 17158 2448 0 _0793_
rlabel metal1 24702 3502 24702 3502 0 _0794_
rlabel metal1 28888 6290 28888 6290 0 _0795_
rlabel metal2 33258 28832 33258 28832 0 _0796_
rlabel metal1 34224 28730 34224 28730 0 _0797_
rlabel metal1 33212 29614 33212 29614 0 _0798_
rlabel metal1 32016 29274 32016 29274 0 _0799_
rlabel metal1 32982 30158 32982 30158 0 _0800_
rlabel metal2 33350 14654 33350 14654 0 _0801_
rlabel metal1 23782 9520 23782 9520 0 _0802_
rlabel metal1 27922 5100 27922 5100 0 _0803_
rlabel metal1 31648 6630 31648 6630 0 _0804_
rlabel metal1 26956 5338 26956 5338 0 _0805_
rlabel metal1 27876 7854 27876 7854 0 _0806_
rlabel metal2 30590 13430 30590 13430 0 _0807_
rlabel metal2 33258 14212 33258 14212 0 _0808_
rlabel metal1 32660 10642 32660 10642 0 _0809_
rlabel metal1 33488 9146 33488 9146 0 _0810_
rlabel metal1 34086 7718 34086 7718 0 _0811_
rlabel metal1 34086 5882 34086 5882 0 _0812_
rlabel metal1 29026 4250 29026 4250 0 _0813_
rlabel metal1 22632 2482 22632 2482 0 _0814_
rlabel metal1 24104 2414 24104 2414 0 _0815_
rlabel metal1 19918 2618 19918 2618 0 _0816_
rlabel metal1 16997 2278 16997 2278 0 _0817_
rlabel metal2 17066 4420 17066 4420 0 _0818_
rlabel metal1 10994 3060 10994 3060 0 _0819_
rlabel metal2 9890 3706 9890 3706 0 _0820_
rlabel metal1 14030 4794 14030 4794 0 _0821_
rlabel metal2 16882 6596 16882 6596 0 _0822_
rlabel metal2 16330 8058 16330 8058 0 _0823_
rlabel metal1 11960 10030 11960 10030 0 _0824_
rlabel metal1 7084 16626 7084 16626 0 _0825_
rlabel metal2 11178 12410 11178 12410 0 _0826_
rlabel metal2 11730 14790 11730 14790 0 _0827_
rlabel metal1 8372 14994 8372 14994 0 _0828_
rlabel metal1 8280 11118 8280 11118 0 _0829_
rlabel metal1 8464 9690 8464 9690 0 _0830_
rlabel metal1 6302 8058 6302 8058 0 _0831_
rlabel metal1 6624 10506 6624 10506 0 _0832_
rlabel metal1 5520 14382 5520 14382 0 _0833_
rlabel metal1 6118 18258 6118 18258 0 _0834_
rlabel metal2 8786 17476 8786 17476 0 _0835_
rlabel metal1 11454 18768 11454 18768 0 _0836_
rlabel metal2 13662 16762 13662 16762 0 _0837_
rlabel metal1 12006 18938 12006 18938 0 _0838_
rlabel metal1 10028 20026 10028 20026 0 _0839_
rlabel metal1 7682 23018 7682 23018 0 _0840_
rlabel metal1 7912 24378 7912 24378 0 _0841_
rlabel metal2 9706 25738 9706 25738 0 _0842_
rlabel metal1 11362 24650 11362 24650 0 _0843_
rlabel metal2 13570 24378 13570 24378 0 _0844_
rlabel metal2 13938 22134 13938 22134 0 _0845_
rlabel metal2 14306 20468 14306 20468 0 _0846_
rlabel metal1 15732 18598 15732 18598 0 _0847_
rlabel metal1 20746 19278 20746 19278 0 _0848_
rlabel metal1 14214 18394 14214 18394 0 _0849_
rlabel metal1 15594 16558 15594 16558 0 _0850_
rlabel metal1 16146 18326 16146 18326 0 _0851_
rlabel metal2 20654 19958 20654 19958 0 _0852_
rlabel metal1 19964 21998 19964 21998 0 _0853_
rlabel metal2 20378 24582 20378 24582 0 _0854_
rlabel metal1 19320 25874 19320 25874 0 _0855_
rlabel metal2 18078 28220 18078 28220 0 _0856_
rlabel metal2 16882 28356 16882 28356 0 _0857_
rlabel metal2 14214 28356 14214 28356 0 _0858_
rlabel metal1 11362 36210 11362 36210 0 _0859_
rlabel metal2 11178 26826 11178 26826 0 _0860_
rlabel metal2 9614 27268 9614 27268 0 _0861_
rlabel metal1 5934 29648 5934 29648 0 _0862_
rlabel metal1 6739 32402 6739 32402 0 _0863_
rlabel metal1 9798 30090 9798 30090 0 _0864_
rlabel metal1 11408 30906 11408 30906 0 _0865_
rlabel metal1 12420 34170 12420 34170 0 _0866_
rlabel metal2 7406 33660 7406 33660 0 _0867_
rlabel metal1 7682 36006 7682 36006 0 _0868_
rlabel metal2 9614 37094 9614 37094 0 _0869_
rlabel metal1 20562 38386 20562 38386 0 _0870_
rlabel metal1 10994 36788 10994 36788 0 _0871_
rlabel metal1 14628 37434 14628 37434 0 _0872_
rlabel metal1 15272 33490 15272 33490 0 _0873_
rlabel metal1 16974 32402 16974 32402 0 _0874_
rlabel metal1 19550 30906 19550 30906 0 _0875_
rlabel metal1 19136 33966 19136 33966 0 _0876_
rlabel metal1 16767 36890 16767 36890 0 _0877_
rlabel metal1 21160 37842 21160 37842 0 _0878_
rlabel metal2 19642 37434 19642 37434 0 _0879_
rlabel metal1 18078 34000 18078 34000 0 _0880_
rlabel metal1 24886 36210 24886 36210 0 _0881_
rlabel metal1 25668 36142 25668 36142 0 _0882_
rlabel metal1 25484 36618 25484 36618 0 _0883_
rlabel metal1 26082 34578 26082 34578 0 _0884_
rlabel metal1 24426 33082 24426 33082 0 _0885_
rlabel metal1 25576 32402 25576 32402 0 _0886_
rlabel metal2 24610 31110 24610 31110 0 _0887_
rlabel metal1 25714 30362 25714 30362 0 _0888_
rlabel metal1 25668 28526 25668 28526 0 _0889_
rlabel metal1 25484 26962 25484 26962 0 _0890_
rlabel metal1 26220 26962 26220 26962 0 _0891_
rlabel metal1 14536 13294 14536 13294 0 _0892_
rlabel metal2 25530 15844 25530 15844 0 _0893_
rlabel metal1 27922 26384 27922 26384 0 _0894_
rlabel metal2 27094 24582 27094 24582 0 _0895_
rlabel metal2 26358 23290 26358 23290 0 _0896_
rlabel metal1 26266 21862 26266 21862 0 _0897_
rlabel metal2 26542 21318 26542 21318 0 _0898_
rlabel metal1 26818 20434 26818 20434 0 _0899_
rlabel metal2 26818 19210 26818 19210 0 _0900_
rlabel metal1 26036 17850 26036 17850 0 _0901_
rlabel metal2 25438 17476 25438 17476 0 _0902_
rlabel metal2 28566 15470 28566 15470 0 _0903_
rlabel metal1 24794 11628 24794 11628 0 _0904_
rlabel metal1 24426 13294 24426 13294 0 _0905_
rlabel metal2 24610 14246 24610 14246 0 _0906_
rlabel metal2 23874 11322 23874 11322 0 _0907_
rlabel metal1 28474 11594 28474 11594 0 _0908_
rlabel metal1 28658 10030 28658 10030 0 _0909_
rlabel metal1 29854 10234 29854 10234 0 _0910_
rlabel metal2 29946 32912 29946 32912 0 _0911_
rlabel metal1 29992 32198 29992 32198 0 _0912_
rlabel metal1 29394 33524 29394 33524 0 _0913_
rlabel metal1 29210 33354 29210 33354 0 _0914_
rlabel metal1 29486 32334 29486 32334 0 _0915_
rlabel via1 29578 32538 29578 32538 0 _0916_
rlabel metal2 29762 31280 29762 31280 0 _0917_
rlabel metal1 28520 30838 28520 30838 0 _0918_
rlabel metal1 28428 31178 28428 31178 0 _0919_
rlabel metal1 28566 31994 28566 31994 0 _0920_
rlabel metal1 28888 32946 28888 32946 0 _0921_
rlabel metal2 27738 37774 27738 37774 0 _0922_
rlabel metal1 28704 37230 28704 37230 0 _0923_
rlabel metal2 28014 37400 28014 37400 0 _0924_
rlabel metal1 28612 37162 28612 37162 0 _0925_
rlabel metal2 28106 36550 28106 36550 0 _0926_
rlabel metal1 28106 35088 28106 35088 0 _0927_
rlabel metal2 28198 35904 28198 35904 0 _0928_
rlabel metal2 28290 35564 28290 35564 0 _0929_
rlabel metal1 28474 35258 28474 35258 0 _0930_
rlabel metal1 28842 35768 28842 35768 0 _0931_
rlabel metal1 28336 34646 28336 34646 0 _0932_
rlabel metal2 28290 34816 28290 34816 0 _0933_
rlabel metal1 27830 35564 27830 35564 0 _0934_
rlabel metal2 28658 35122 28658 35122 0 _0935_
rlabel metal1 29072 32878 29072 32878 0 _0936_
rlabel metal1 27784 34170 27784 34170 0 _0937_
rlabel metal1 28566 35666 28566 35666 0 _0938_
rlabel metal1 28428 32946 28428 32946 0 _0939_
rlabel metal1 28612 32742 28612 32742 0 _0940_
rlabel metal1 28934 31926 28934 31926 0 _0941_
rlabel metal1 29946 31824 29946 31824 0 _0942_
rlabel metal1 30452 31790 30452 31790 0 _0943_
rlabel metal2 31786 28356 31786 28356 0 _0944_
rlabel metal1 32476 28118 32476 28118 0 _0945_
rlabel metal2 32338 23936 32338 23936 0 _0946_
rlabel metal1 33074 22542 33074 22542 0 _0947_
rlabel metal1 29578 21590 29578 21590 0 _0948_
rlabel metal2 30682 22848 30682 22848 0 _0949_
rlabel metal1 29762 21998 29762 21998 0 _0950_
rlabel metal2 32890 21794 32890 21794 0 _0951_
rlabel metal1 32292 22202 32292 22202 0 _0952_
rlabel metal1 32246 22678 32246 22678 0 _0953_
rlabel metal2 33994 26554 33994 26554 0 _0954_
rlabel metal2 36478 27132 36478 27132 0 _0955_
rlabel metal1 32522 25908 32522 25908 0 _0956_
rlabel metal1 33994 28118 33994 28118 0 _0957_
rlabel metal1 32522 28424 32522 28424 0 _0958_
rlabel metal1 30452 28050 30452 28050 0 _0959_
rlabel metal1 36662 27030 36662 27030 0 _0960_
rlabel metal2 32614 25670 32614 25670 0 _0961_
rlabel metal1 33166 22610 33166 22610 0 _0962_
rlabel metal2 33534 24208 33534 24208 0 _0963_
rlabel metal2 33258 24514 33258 24514 0 _0964_
rlabel metal1 32522 22542 32522 22542 0 _0965_
rlabel metal2 33810 23834 33810 23834 0 _0966_
rlabel via1 32811 22678 32811 22678 0 _0967_
rlabel metal1 30038 22032 30038 22032 0 _0968_
rlabel metal2 29394 21692 29394 21692 0 _0969_
rlabel metal2 28750 21590 28750 21590 0 _0970_
rlabel metal2 29210 21216 29210 21216 0 _0971_
rlabel metal2 28750 15980 28750 15980 0 _0972_
rlabel metal1 29578 15028 29578 15028 0 _0973_
rlabel metal1 30360 14450 30360 14450 0 _0974_
rlabel metal2 29854 15164 29854 15164 0 _0975_
rlabel metal1 29394 15130 29394 15130 0 _0976_
rlabel metal1 28796 17170 28796 17170 0 _0977_
rlabel metal2 28842 18462 28842 18462 0 _0978_
rlabel metal2 28658 18054 28658 18054 0 _0979_
rlabel metal1 29716 17306 29716 17306 0 _0980_
rlabel metal1 28428 17306 28428 17306 0 _0981_
rlabel metal2 29486 17068 29486 17068 0 _0982_
rlabel metal2 30038 16388 30038 16388 0 _0983_
rlabel metal1 28842 13872 28842 13872 0 _0984_
rlabel metal1 32867 15946 32867 15946 0 _0985_
rlabel metal1 28198 15674 28198 15674 0 _0986_
rlabel metal2 27738 15334 27738 15334 0 _0987_
rlabel metal2 29026 14892 29026 14892 0 _0988_
rlabel metal2 29118 14076 29118 14076 0 _0989_
rlabel metal1 28888 13770 28888 13770 0 _0990_
rlabel metal1 28336 14586 28336 14586 0 _0991_
rlabel metal2 26266 1962 26266 1962 0 clk_in
rlabel metal2 21850 33184 21850 33184 0 clknet_0_clk_in
rlabel metal1 33258 22678 33258 22678 0 clknet_0_ref_in
rlabel metal2 33626 35598 33626 35598 0 clknet_0_vco_in
rlabel metal2 34362 20672 34362 20672 0 clknet_1_0__leaf_ref_in
rlabel metal2 32798 32368 32798 32368 0 clknet_1_0__leaf_vco_in
rlabel metal1 36478 25738 36478 25738 0 clknet_1_1__leaf_ref_in
rlabel metal2 34086 37298 34086 37298 0 clknet_1_1__leaf_vco_in
rlabel metal1 12282 2958 12282 2958 0 clknet_4_0_0_clk_in
rlabel metal1 6578 28118 6578 28118 0 clknet_4_10_0_clk_in
rlabel metal1 12006 37094 12006 37094 0 clknet_4_11_0_clk_in
rlabel metal1 20102 22066 20102 22066 0 clknet_4_12_0_clk_in
rlabel metal1 22034 24650 22034 24650 0 clknet_4_13_0_clk_in
rlabel metal2 16882 37434 16882 37434 0 clknet_4_14_0_clk_in
rlabel metal1 22034 33524 22034 33524 0 clknet_4_15_0_clk_in
rlabel metal1 17158 3978 17158 3978 0 clknet_4_1_0_clk_in
rlabel metal1 6348 12818 6348 12818 0 clknet_4_2_0_clk_in
rlabel metal1 6440 15538 6440 15538 0 clknet_4_3_0_clk_in
rlabel metal2 22034 3808 22034 3808 0 clknet_4_4_0_clk_in
rlabel metal2 29762 4284 29762 4284 0 clknet_4_5_0_clk_in
rlabel metal1 21620 12274 21620 12274 0 clknet_4_6_0_clk_in
rlabel metal1 24932 12274 24932 12274 0 clknet_4_7_0_clk_in
rlabel metal1 6670 22644 6670 22644 0 clknet_4_8_0_clk_in
rlabel metal2 11178 24786 11178 24786 0 clknet_4_9_0_clk_in
rlabel metal2 36938 38607 36938 38607 0 corner[0]
rlabel metal2 37122 34969 37122 34969 0 corner[1]
rlabel metal2 37122 31501 37122 31501 0 corner[2]
rlabel metal1 26726 19482 26726 19482 0 d2.r_reg\[10\]
rlabel metal2 25622 20672 25622 20672 0 d2.r_reg\[11\]
rlabel metal1 25668 21930 25668 21930 0 d2.r_reg\[12\]
rlabel metal1 25760 23086 25760 23086 0 d2.r_reg\[13\]
rlabel metal1 25438 24922 25438 24922 0 d2.r_reg\[14\]
rlabel metal2 26082 26112 26082 26112 0 d2.r_reg\[15\]
rlabel metal1 24840 25874 24840 25874 0 d2.r_reg\[16\]
rlabel metal2 22678 26928 22678 26928 0 d2.r_reg\[17\]
rlabel metal1 24242 28526 24242 28526 0 d2.r_reg\[18\]
rlabel metal2 23598 29886 23598 29886 0 d2.r_reg\[19\]
rlabel metal2 25990 10370 25990 10370 0 d2.r_reg\[1\]
rlabel metal2 23874 30430 23874 30430 0 d2.r_reg\[20\]
rlabel metal1 24242 32538 24242 32538 0 d2.r_reg\[21\]
rlabel metal1 24334 32878 24334 32878 0 d2.r_reg\[22\]
rlabel metal2 23966 34816 23966 34816 0 d2.r_reg\[23\]
rlabel metal1 25760 36754 25760 36754 0 d2.r_reg\[24\]
rlabel metal1 23690 36550 23690 36550 0 d2.r_reg\[25\]
rlabel metal2 19918 35428 19918 35428 0 d2.r_reg\[26\]
rlabel metal1 20148 36142 20148 36142 0 d2.r_reg\[27\]
rlabel metal1 20378 38250 20378 38250 0 d2.r_reg\[28\]
rlabel metal1 18446 36142 18446 36142 0 d2.r_reg\[29\]
rlabel metal2 25622 10642 25622 10642 0 d2.r_reg\[2\]
rlabel metal1 18768 33626 18768 33626 0 d2.r_reg\[30\]
rlabel metal1 19412 31858 19412 31858 0 d2.r_reg\[31\]
rlabel metal1 17342 30328 17342 30328 0 d2.r_reg\[32\]
rlabel metal1 15594 32742 15594 32742 0 d2.r_reg\[33\]
rlabel metal1 15226 37094 15226 37094 0 d2.r_reg\[34\]
rlabel metal2 13110 36414 13110 36414 0 d2.r_reg\[35\]
rlabel metal1 12558 36040 12558 36040 0 d2.r_reg\[36\]
rlabel metal1 10856 35462 10856 35462 0 d2.r_reg\[37\]
rlabel metal1 9568 34034 9568 34034 0 d2.r_reg\[38\]
rlabel metal2 12190 33320 12190 33320 0 d2.r_reg\[39\]
rlabel metal2 24702 11356 24702 11356 0 d2.r_reg\[3\]
rlabel metal2 11546 32334 11546 32334 0 d2.r_reg\[40\]
rlabel metal1 11500 30226 11500 30226 0 d2.r_reg\[41\]
rlabel metal1 8878 30362 8878 30362 0 d2.r_reg\[42\]
rlabel metal2 8326 29954 8326 29954 0 d2.r_reg\[43\]
rlabel metal1 9200 27098 9200 27098 0 d2.r_reg\[44\]
rlabel metal1 11224 28186 11224 28186 0 d2.r_reg\[45\]
rlabel metal1 14674 28084 14674 28084 0 d2.r_reg\[46\]
rlabel metal1 16560 28118 16560 28118 0 d2.r_reg\[47\]
rlabel metal1 18538 28594 18538 28594 0 d2.r_reg\[48\]
rlabel metal1 19228 26418 19228 26418 0 d2.r_reg\[49\]
rlabel metal1 22908 12410 22908 12410 0 d2.r_reg\[4\]
rlabel metal1 19504 24786 19504 24786 0 d2.r_reg\[50\]
rlabel metal1 18883 21998 18883 21998 0 d2.r_reg\[51\]
rlabel metal2 21114 20468 21114 20468 0 d2.r_reg\[52\]
rlabel metal2 20746 17510 20746 17510 0 d2.r_reg\[53\]
rlabel metal1 17434 17238 17434 17238 0 d2.r_reg\[54\]
rlabel metal1 15180 17714 15180 17714 0 d2.r_reg\[55\]
rlabel metal1 14628 19754 14628 19754 0 d2.r_reg\[56\]
rlabel metal2 13478 21012 13478 21012 0 d2.r_reg\[57\]
rlabel metal1 13064 21998 13064 21998 0 d2.r_reg\[58\]
rlabel metal2 12190 24276 12190 24276 0 d2.r_reg\[59\]
rlabel metal1 23828 12818 23828 12818 0 d2.r_reg\[5\]
rlabel metal2 9706 23188 9706 23188 0 d2.r_reg\[60\]
rlabel metal1 8280 24242 8280 24242 0 d2.r_reg\[61\]
rlabel metal1 8924 23086 8924 23086 0 d2.r_reg\[62\]
rlabel metal1 9798 19312 9798 19312 0 d2.r_reg\[63\]
rlabel metal2 11638 19278 11638 19278 0 d2.r_reg\[64\]
rlabel metal2 13018 15878 13018 15878 0 d2.r_reg\[65\]
rlabel metal1 10902 16456 10902 16456 0 d2.r_reg\[66\]
rlabel metal2 6854 16796 6854 16796 0 d2.r_reg\[67\]
rlabel metal1 8004 15674 8004 15674 0 d2.r_reg\[68\]
rlabel metal2 7038 11118 7038 11118 0 d2.r_reg\[69\]
rlabel metal1 24610 16150 24610 16150 0 d2.r_reg\[6\]
rlabel metal1 7038 8806 7038 8806 0 d2.r_reg\[70\]
rlabel metal2 8234 9214 8234 9214 0 d2.r_reg\[71\]
rlabel metal1 9614 11866 9614 11866 0 d2.r_reg\[72\]
rlabel metal2 10074 14688 10074 14688 0 d2.r_reg\[73\]
rlabel metal2 12190 14178 12190 14178 0 d2.r_reg\[74\]
rlabel metal1 10994 11866 10994 11866 0 d2.r_reg\[75\]
rlabel metal2 12742 10540 12742 10540 0 d2.r_reg\[76\]
rlabel metal1 14582 8500 14582 8500 0 d2.r_reg\[77\]
rlabel metal2 15778 6018 15778 6018 0 d2.r_reg\[78\]
rlabel metal1 14720 6426 14720 6426 0 d2.r_reg\[79\]
rlabel metal1 24840 17034 24840 17034 0 d2.r_reg\[7\]
rlabel metal2 12650 4182 12650 4182 0 d2.r_reg\[80\]
rlabel metal1 12512 4114 12512 4114 0 d2.r_reg\[81\]
rlabel metal2 14582 4284 14582 4284 0 d2.r_reg\[82\]
rlabel metal2 18906 4352 18906 4352 0 d2.r_reg\[83\]
rlabel metal1 20332 3026 20332 3026 0 d2.r_reg\[84\]
rlabel metal1 23368 4046 23368 4046 0 d2.r_reg\[85\]
rlabel metal1 28566 4454 28566 4454 0 d2.r_reg\[86\]
rlabel metal1 31188 5270 31188 5270 0 d2.r_reg\[87\]
rlabel metal1 32660 6766 32660 6766 0 d2.r_reg\[88\]
rlabel metal1 33258 8874 33258 8874 0 d2.r_reg\[89\]
rlabel metal2 23690 17884 23690 17884 0 d2.r_reg\[8\]
rlabel metal1 33718 11254 33718 11254 0 d2.r_reg\[90\]
rlabel metal2 33166 12279 33166 12279 0 d2.r_reg\[91\]
rlabel metal2 30038 11968 30038 11968 0 d2.r_reg\[92\]
rlabel metal1 30590 8602 30590 8602 0 d2.r_reg\[93\]
rlabel metal2 27646 5780 27646 5780 0 d2.r_reg\[94\]
rlabel metal1 30636 6698 30636 6698 0 d2.r_reg\[95\]
rlabel metal2 25070 19550 25070 19550 0 d2.r_reg\[9\]
rlabel metal1 28796 10574 28796 10574 0 d2.t_load\[0\]
rlabel metal1 27876 20570 27876 20570 0 d2.t_load\[10\]
rlabel metal1 28106 21658 28106 21658 0 d2.t_load\[11\]
rlabel metal2 28014 30192 28014 30192 0 d2.t_load\[12\]
rlabel metal1 28566 29614 28566 29614 0 d2.t_load\[13\]
rlabel metal2 28382 26163 28382 26163 0 d2.t_load\[14\]
rlabel metal1 26312 26214 26312 26214 0 d2.t_load\[15\]
rlabel metal1 24886 28050 24886 28050 0 d2.t_load\[16\]
rlabel metal1 24702 27030 24702 27030 0 d2.t_load\[17\]
rlabel metal1 28842 28560 28842 28560 0 d2.t_load\[18\]
rlabel metal1 24518 30226 24518 30226 0 d2.t_load\[19\]
rlabel metal1 27646 12274 27646 12274 0 d2.t_load\[1\]
rlabel metal1 24426 32266 24426 32266 0 d2.t_load\[20\]
rlabel metal1 27186 31858 27186 31858 0 d2.t_load\[21\]
rlabel metal2 24978 33728 24978 33728 0 d2.t_load\[22\]
rlabel metal1 25622 35054 25622 35054 0 d2.t_load\[23\]
rlabel metal1 25346 36822 25346 36822 0 d2.t_load\[24\]
rlabel metal1 28750 36074 28750 36074 0 d2.t_load\[25\]
rlabel metal2 20010 35943 20010 35943 0 d2.t_load\[26\]
rlabel metal1 21068 37910 21068 37910 0 d2.t_load\[27\]
rlabel metal1 20286 38318 20286 38318 0 d2.t_load\[28\]
rlabel metal1 18078 37094 18078 37094 0 d2.t_load\[29\]
rlabel metal2 26634 11492 26634 11492 0 d2.t_load\[2\]
rlabel metal1 19734 32538 19734 32538 0 d2.t_load\[30\]
rlabel metal1 19504 30702 19504 30702 0 d2.t_load\[31\]
rlabel metal2 16054 31518 16054 31518 0 d2.t_load\[32\]
rlabel metal1 17756 32742 17756 32742 0 d2.t_load\[33\]
rlabel metal1 14674 37230 14674 37230 0 d2.t_load\[34\]
rlabel metal2 13478 37638 13478 37638 0 d2.t_load\[35\]
rlabel metal1 10258 36720 10258 36720 0 d2.t_load\[36\]
rlabel metal1 8188 36006 8188 36006 0 d2.t_load\[37\]
rlabel metal2 8510 33490 8510 33490 0 d2.t_load\[38\]
rlabel metal1 12972 33830 12972 33830 0 d2.t_load\[39\]
rlabel metal1 25070 12308 25070 12308 0 d2.t_load\[3\]
rlabel metal2 12190 31518 12190 31518 0 d2.t_load\[40\]
rlabel metal1 10166 30294 10166 30294 0 d2.t_load\[41\]
rlabel metal2 8234 31280 8234 31280 0 d2.t_load\[42\]
rlabel metal1 8970 28934 8970 28934 0 d2.t_load\[43\]
rlabel metal1 13570 37774 13570 37774 0 d2.t_load\[44\]
rlabel metal1 14260 26418 14260 26418 0 d2.t_load\[45\]
rlabel metal1 15870 27948 15870 27948 0 d2.t_load\[46\]
rlabel metal2 17618 26826 17618 26826 0 d2.t_load\[47\]
rlabel metal2 18446 27948 18446 27948 0 d2.t_load\[48\]
rlabel metal2 19918 25772 19918 25772 0 d2.t_load\[49\]
rlabel metal1 27048 13838 27048 13838 0 d2.t_load\[4\]
rlabel metal1 19964 23154 19964 23154 0 d2.t_load\[50\]
rlabel metal1 20746 21658 20746 21658 0 d2.t_load\[51\]
rlabel metal2 20838 18938 20838 18938 0 d2.t_load\[52\]
rlabel metal2 19458 19754 19458 19754 0 d2.t_load\[53\]
rlabel metal1 17388 18734 17388 18734 0 d2.t_load\[54\]
rlabel metal1 16882 19210 16882 19210 0 d2.t_load\[55\]
rlabel metal2 14306 36861 14306 36861 0 d2.t_load\[56\]
rlabel metal1 14812 21590 14812 21590 0 d2.t_load\[57\]
rlabel metal1 11178 23766 11178 23766 0 d2.t_load\[58\]
rlabel metal2 12098 25194 12098 25194 0 d2.t_load\[59\]
rlabel metal2 26726 14144 26726 14144 0 d2.t_load\[5\]
rlabel metal1 10764 25738 10764 25738 0 d2.t_load\[60\]
rlabel metal2 9246 23766 9246 23766 0 d2.t_load\[61\]
rlabel metal1 8786 23664 8786 23664 0 d2.t_load\[62\]
rlabel metal2 11546 20230 11546 20230 0 d2.t_load\[63\]
rlabel metal2 12190 17578 12190 17578 0 d2.t_load\[64\]
rlabel metal1 16514 16014 16514 16014 0 d2.t_load\[65\]
rlabel metal2 25622 14960 25622 14960 0 d2.t_load\[6\]
rlabel metal1 25254 17170 25254 17170 0 d2.t_load\[7\]
rlabel metal1 25484 17578 25484 17578 0 d2.t_load\[8\]
rlabel metal1 28244 8602 28244 8602 0 d2.t_load\[93\]
rlabel metal1 28382 5882 28382 5882 0 d2.t_load\[94\]
rlabel metal2 31326 6494 31326 6494 0 d2.t_load\[95\]
rlabel metal1 26082 19278 26082 19278 0 d2.t_load\[9\]
rlabel metal1 33120 29274 33120 29274 0 d5.fll_core.corner_tmp\[0\]
rlabel metal2 33994 30124 33994 30124 0 d5.fll_core.corner_tmp\[1\]
rlabel metal1 31510 29274 31510 29274 0 d5.fll_core.corner_tmp\[2\]
rlabel metal1 32131 32402 32131 32402 0 d5.fll_core.counter1.count\[0\]
rlabel metal1 30912 31790 30912 31790 0 d5.fll_core.counter1.count\[1\]
rlabel metal1 31372 32402 31372 32402 0 d5.fll_core.counter1.count\[2\]
rlabel metal2 27738 32708 27738 32708 0 d5.fll_core.counter1.count\[3\]
rlabel metal1 31050 34578 31050 34578 0 d5.fll_core.counter1.count\[4\]
rlabel metal1 29440 35734 29440 35734 0 d5.fll_core.counter1.count\[5\]
rlabel metal1 30912 34918 30912 34918 0 d5.fll_core.counter1.count\[6\]
rlabel metal1 30590 36754 30590 36754 0 d5.fll_core.counter1.count\[7\]
rlabel metal1 28428 38318 28428 38318 0 d5.fll_core.counter1.count\[8\]
rlabel metal2 29854 36924 29854 36924 0 d5.fll_core.counter1.count\[9\]
rlabel metal2 34086 17374 34086 17374 0 d5.fll_core.counter2.count\[0\]
rlabel metal1 33120 17714 33120 17714 0 d5.fll_core.counter2.count\[1\]
rlabel metal1 35144 17578 35144 17578 0 d5.fll_core.counter2.count\[2\]
rlabel metal2 35650 14654 35650 14654 0 d5.fll_core.counter2.count\[3\]
rlabel metal2 36294 15164 36294 15164 0 d5.fll_core.counter2.count\[4\]
rlabel metal1 32568 15674 32568 15674 0 d5.fll_core.counter2.count\[5\]
rlabel metal1 30774 14892 30774 14892 0 d5.fll_core.counter2.count\[6\]
rlabel metal1 32108 16966 32108 16966 0 d5.fll_core.counter2.count\[7\]
rlabel metal1 32062 18394 32062 18394 0 d5.fll_core.counter2.count\[8\]
rlabel metal2 31878 18938 31878 18938 0 d5.fll_core.counter2.count\[9\]
rlabel metal1 32246 30226 32246 30226 0 d5.fll_core.counter_reset
rlabel metal1 18814 20910 18814 20910 0 d5.fll_core.strobe
rlabel metal1 33534 28084 33534 28084 0 d5.fll_core.tmp\[0\]
rlabel metal1 33350 26996 33350 26996 0 d5.fll_core.tmp\[1\]
rlabel metal2 36662 27676 36662 27676 0 d5.fll_core.tmp\[2\]
rlabel metal1 32384 25194 32384 25194 0 d5.fll_core.tmp\[3\]
rlabel metal2 32522 23426 32522 23426 0 d5.fll_core.tmp\[4\]
rlabel metal2 36846 23970 36846 23970 0 d5.fll_core.tmp\[5\]
rlabel metal1 33580 23290 33580 23290 0 d5.fll_core.tmp\[6\]
rlabel metal2 33626 22610 33626 22610 0 d5.fll_core.tmp\[7\]
rlabel metal1 19642 20366 19642 20366 0 d5.fll_core.tmp\[8\]
rlabel metal1 18124 19482 18124 19482 0 d5.fll_core.tmp\[9\]
rlabel metal2 14582 25500 14582 25500 0 d5.mux01.out\[0\]
rlabel metal2 14214 26622 14214 26622 0 d5.mux01.out\[1\]
rlabel metal2 18354 26248 18354 26248 0 d5.mux01.out\[2\]
rlabel metal1 16606 25330 16606 25330 0 d5.mux01.out\[3\]
rlabel metal2 17158 24412 17158 24412 0 d5.mux01.out\[4\]
rlabel metal1 15686 23154 15686 23154 0 d5.mux01.out\[5\]
rlabel metal1 17342 22542 17342 22542 0 d5.mux01.out\[6\]
rlabel metal1 17250 20570 17250 20570 0 d5.mux01.out\[7\]
rlabel metal1 19412 19278 19412 19278 0 d5.mux01.out\[8\]
rlabel metal1 16238 19754 16238 19754 0 d5.mux01.out\[9\]
rlabel metal2 1794 39355 1794 39355 0 dac[0]
rlabel metal2 4738 39355 4738 39355 0 dac[1]
rlabel metal2 7682 39355 7682 39355 0 dac[2]
rlabel metal1 10212 38522 10212 38522 0 dac[3]
rlabel metal1 12144 38522 12144 38522 0 dac[4]
rlabel metal2 16330 39355 16330 39355 0 dac[5]
rlabel metal2 19274 38250 19274 38250 0 dac[6]
rlabel metal1 22356 38522 22356 38522 0 dac[7]
rlabel metal2 31786 1588 31786 1588 0 load
rlabel metal1 25530 10642 25530 10642 0 net1
rlabel metal2 8142 38148 8142 38148 0 net10
rlabel metal2 10166 38148 10166 38148 0 net11
rlabel metal1 10764 38318 10764 38318 0 net12
rlabel metal2 15778 38148 15778 38148 0 net13
rlabel metal2 19090 38148 19090 38148 0 net14
rlabel metal2 14766 37570 14766 37570 0 net15
rlabel metal1 36317 2414 36317 2414 0 net16
rlabel metal1 1932 35054 1932 35054 0 net17
rlabel metal2 1794 28390 1794 28390 0 net18
rlabel metal1 1886 31790 1886 31790 0 net19
rlabel metal1 25369 2346 25369 2346 0 net2
rlabel metal1 4830 3026 4830 3026 0 net20
rlabel metal1 4416 5678 4416 5678 0 net21
rlabel metal1 1794 9588 1794 9588 0 net22
rlabel metal1 1794 13260 1794 13260 0 net23
rlabel metal1 1794 17238 1794 17238 0 net24
rlabel metal1 1978 20434 1978 20434 0 net25
rlabel metal1 2024 24174 2024 24174 0 net26
rlabel metal1 1840 28050 1840 28050 0 net27
rlabel metal1 20056 8330 20056 8330 0 net28
rlabel metal2 17618 4046 17618 4046 0 net29
rlabel metal2 25254 2720 25254 2720 0 net3
rlabel metal1 12880 5134 12880 5134 0 net30
rlabel metal1 10810 4148 10810 4148 0 net31
rlabel metal1 13064 3366 13064 3366 0 net32
rlabel metal1 16675 3434 16675 3434 0 net33
rlabel metal2 4462 2176 4462 2176 0 net34
rlabel metal2 1794 2244 1794 2244 0 net35
rlabel metal1 24702 3978 24702 3978 0 net36
rlabel metal2 36938 5202 36938 5202 0 net37
rlabel metal2 33534 6188 33534 6188 0 net38
rlabel metal1 34178 8602 34178 8602 0 net39
rlabel metal1 34868 2618 34868 2618 0 net4
rlabel metal1 36409 9486 36409 9486 0 net40
rlabel metal2 33258 11968 33258 11968 0 net41
rlabel metal1 33304 12342 33304 12342 0 net42
rlabel metal1 36984 27438 36984 27438 0 net43
rlabel metal1 25576 38522 25576 38522 0 net44
rlabel metal1 29394 38454 29394 38454 0 net45
rlabel metal1 34132 38522 34132 38522 0 net46
rlabel metal2 34730 38148 34730 38148 0 net5
rlabel metal1 35788 31450 35788 31450 0 net6
rlabel metal1 34178 31450 34178 31450 0 net7
rlabel metal1 1978 38352 1978 38352 0 net8
rlabel metal1 4968 37978 4968 37978 0 net9
rlabel metal2 29026 1554 29026 1554 0 read
rlabel metal1 35696 22678 35696 22678 0 ref_in
rlabel metal2 23506 1622 23506 1622 0 reset
rlabel metal2 34546 1588 34546 1588 0 s_in
rlabel metal2 37306 1520 37306 1520 0 s_out
rlabel metal3 1142 35020 1142 35020 0 slope_ctrl[0]
rlabel metal2 1610 38335 1610 38335 0 slope_ctrl[1]
rlabel metal3 1142 31348 1142 31348 0 slope_ctrl[2]
rlabel metal3 1142 1972 1142 1972 0 vbias1[0]
rlabel metal3 1142 5644 1142 5644 0 vbias1[1]
rlabel metal3 1142 9316 1142 9316 0 vbias1[2]
rlabel metal3 1142 12988 1142 12988 0 vbias1[3]
rlabel metal3 1142 16660 1142 16660 0 vbias1[4]
rlabel metal3 1142 20332 1142 20332 0 vbias1[5]
rlabel metal3 1142 24004 1142 24004 0 vbias1[6]
rlabel metal3 1142 27676 1142 27676 0 vbias1[7]
rlabel metal2 20746 1520 20746 1520 0 vbias2[0]
rlabel metal2 17986 1520 17986 1520 0 vbias2[1]
rlabel metal2 15226 1095 15226 1095 0 vbias2[2]
rlabel metal2 12466 1690 12466 1690 0 vbias2[3]
rlabel metal2 9706 1520 9706 1520 0 vbias2[4]
rlabel metal2 6946 1520 6946 1520 0 vbias2[5]
rlabel metal2 4186 1520 4186 1520 0 vbias2[6]
rlabel metal2 1426 1520 1426 1520 0 vbias2[7]
rlabel metal2 36938 2397 36938 2397 0 vbias3[0]
rlabel metal2 37122 5593 37122 5593 0 vbias3[1]
rlabel via2 36938 9333 36938 9333 0 vbias3[2]
rlabel metal2 37122 13073 37122 13073 0 vbias3[3]
rlabel metal2 37122 16541 37122 16541 0 vbias3[4]
rlabel via2 36938 20315 36938 20315 0 vbias3[5]
rlabel via2 37122 24021 37122 24021 0 vbias3[6]
rlabel metal2 37122 27625 37122 27625 0 vbias3[7]
rlabel metal2 31142 37410 31142 37410 0 vco_in
<< properties >>
string FIXED_BBOX 0 0 38749 40893
<< end >>
