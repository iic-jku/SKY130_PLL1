magic
tech sky130A
magscale 1 2
timestamp 1668357910
<< locali >>
rect 108 306 142 455
rect 1068 306 1102 455
rect 300 -543 334 -403
rect 876 -543 910 -403
<< metal1 >>
rect 584 -32 626 85
rect -42 -74 626 -32
rect 584 -191 626 -74
<< metal2 >>
rect 584 -32 626 166
rect 584 -74 1252 -32
rect 584 -263 626 -74
use sinv2_n  sinv2_n_0
timestamp 1668357910
transform 1 0 605 0 1 -333
box -455 -280 455 280
use sinv2_p  sinv2_p_0
timestamp 1668357910
transform 1 0 605 0 1 236
box -647 -289 647 289
<< end >>
