magic
tech sky130A
magscale 1 2
timestamp 1668357910
<< metal1 >>
rect 807 1886 871 1892
rect -139 1822 807 1886
rect -139 1463 -75 1822
rect 807 1816 871 1822
rect 1476 1719 1543 1876
rect -139 1393 -75 1399
rect -42 1677 1543 1719
rect -42 581 0 1677
rect 428 1571 483 1577
rect 422 1516 428 1571
rect 483 1516 920 1571
rect 1476 1520 1543 1677
rect 1788 1672 1794 1724
rect 1846 1672 1852 1724
rect 428 1510 483 1516
rect 2730 1407 2788 1413
rect -42 539 147 581
rect 878 534 884 586
rect 936 534 942 586
rect 1788 534 1794 586
rect 1846 534 1852 586
rect 2730 269 2788 1349
rect 2730 205 2788 211
<< via1 >>
rect 807 1822 871 1886
rect -139 1399 -75 1463
rect 428 1516 483 1571
rect 1794 1672 1846 1724
rect 2730 1349 2788 1407
rect 884 534 936 586
rect 1794 534 1846 586
rect 2730 211 2788 269
<< metal2 >>
rect 772 1987 1050 2057
rect 427 1571 485 1929
rect 801 1822 807 1886
rect 871 1822 877 1886
rect -139 1516 428 1571
rect 483 1516 489 1571
rect -139 1513 483 1516
rect -145 1399 -139 1463
rect -75 1399 -69 1463
rect -139 269 -75 1399
rect 80 919 138 1513
rect 428 1510 483 1513
rect 810 1488 868 1822
rect 1337 1719 1395 1917
rect 1794 1724 1846 1730
rect 1337 1677 1794 1719
rect 1528 1488 1586 1677
rect 1794 1666 1846 1672
rect 1060 1348 1337 1418
rect 1900 919 1958 2057
rect 2592 1999 2794 2057
rect 2730 1677 2772 1719
rect 2496 1349 2730 1407
rect 2788 1349 2794 1407
rect 80 861 147 919
rect 772 849 1048 919
rect 1682 849 1958 919
rect 884 586 936 592
rect 878 539 884 581
rect 1794 586 1846 592
rect 1788 539 1794 581
rect 884 528 936 534
rect 2730 539 2772 581
rect 1794 528 1846 534
rect -139 211 234 269
rect 676 211 1144 281
rect 1586 211 2054 281
rect 2496 211 2730 269
rect 2788 211 2794 269
use diff_n  diff_n_0
timestamp 1668357910
transform 1 0 1557 0 1 1418
box -359 -280 359 280
use diff_p  diff_p_0
timestamp 1668357910
transform 1 0 1366 0 1 1987
box -455 -289 455 289
use inv_simple1  inv_simple1_0
timestamp 1668357910
transform 1 0 53 0 1 613
box -53 -613 858 525
use inv_simple1  inv_simple1_1
timestamp 1668357910
transform 1 0 963 0 1 613
box -53 -613 858 525
use inv_simple1  inv_simple1_2
timestamp 1668357910
transform 1 0 1873 0 1 613
box -53 -613 858 525
use inv_simple1  inv_simple1_3
timestamp 1668357910
transform 1 0 1873 0 1 1751
box -53 -613 858 525
use diff_n  sky130_fd_pr__nfet_01v8_2AA63J_0
timestamp 1668357910
transform 1 0 839 0 1 1418
box -359 -280 359 280
use diff_p  sky130_fd_pr__pfet_01v8_X6FFBL_0
timestamp 1668357910
transform 1 0 456 0 1 1987
box -455 -289 455 289
<< labels >>
rlabel metal2 2730 539 2772 581 0 nclk
port 1 n
rlabel metal2 2730 1677 2772 1719 0 clk
port 2 n
rlabel metal2 2736 1999 2794 2057 5 vdd
port 4 n
rlabel metal1 -42 1677 0 1719 6 clk_in
port 5 n
rlabel metal1 -139 1822 -75 1886 7 vss
port 3 n
<< end >>
