magic
tech sky130A
magscale 1 2
timestamp 1668153059
<< pwell >>
rect 1435 -70 1821 0
rect 3455 -70 3841 0
rect 1435 -256 2087 -70
rect 3189 -256 3841 -70
<< metal1 >>
rect 609 381 615 443
rect 677 381 710 443
rect 772 381 807 443
rect 869 381 903 443
rect 965 381 999 443
rect 1061 381 1095 443
rect 1157 381 1191 443
rect 1253 381 1287 443
rect 1349 381 1383 443
rect 1445 381 1481 443
rect 1543 381 1549 443
rect 671 350 717 381
rect 863 350 909 381
rect 1055 350 1101 381
rect 1247 350 1293 381
rect 1439 350 1485 381
rect 2226 350 2272 740
rect 3004 350 3050 728
rect 3330 565 3382 571
rect 3330 507 3382 513
rect 3333 359 3378 507
rect 3730 381 3736 443
rect 3798 381 3831 443
rect 3893 381 3928 443
rect 3990 381 4024 443
rect 4086 381 4120 443
rect 4182 381 4216 443
rect 4278 381 4312 443
rect 4374 381 4408 443
rect 4470 381 4504 443
rect 4566 381 4602 443
rect 4664 381 4670 443
rect 3330 353 3382 359
rect 3330 295 3382 301
rect 3786 343 3842 350
rect 3786 287 3788 343
rect 3841 287 3842 343
rect 3786 280 3842 287
rect 3978 343 4034 350
rect 3978 287 3980 343
rect 4033 287 4034 343
rect 3978 280 4034 287
rect 4170 343 4226 350
rect 4170 287 4172 343
rect 4225 287 4226 343
rect 4170 280 4226 287
rect 4362 343 4418 350
rect 4362 287 4364 343
rect 4417 287 4418 343
rect 4362 280 4418 287
rect 4554 343 4611 350
rect 4554 287 4556 343
rect 4609 287 4611 343
rect 4554 280 4611 287
rect 2168 132 2330 178
rect 2946 132 3108 178
rect 2365 -248 2911 -202
<< via1 >>
rect 615 381 677 443
rect 710 381 772 443
rect 807 381 869 443
rect 903 381 965 443
rect 999 381 1061 443
rect 1095 381 1157 443
rect 1191 381 1253 443
rect 1287 381 1349 443
rect 1383 381 1445 443
rect 1481 381 1543 443
rect 3330 513 3382 565
rect 3736 381 3798 443
rect 3831 381 3893 443
rect 3928 381 3990 443
rect 4024 381 4086 443
rect 4120 381 4182 443
rect 4216 381 4278 443
rect 4312 381 4374 443
rect 4408 381 4470 443
rect 4504 381 4566 443
rect 4602 381 4664 443
rect 3330 301 3382 353
rect 3788 287 3841 343
rect 3980 287 4033 343
rect 4172 287 4225 343
rect 4364 287 4417 343
rect 4556 287 4609 343
<< metal2 >>
rect 0 849 139 919
rect 2499 849 2777 919
rect 5137 849 5276 919
rect 1192 443 1254 821
rect 3333 565 3378 779
rect 3324 513 3330 565
rect 3382 513 3388 565
rect 609 381 615 443
rect 677 381 710 443
rect 772 381 807 443
rect 869 381 903 443
rect 965 381 999 443
rect 1061 381 1095 443
rect 1157 381 1191 443
rect 1253 381 1287 443
rect 1349 381 1383 443
rect 1445 381 1481 443
rect 1543 381 3736 443
rect 3798 381 3831 443
rect 3893 381 3928 443
rect 3990 381 4024 443
rect 4086 381 4120 443
rect 4182 381 4216 443
rect 4278 381 4312 443
rect 4374 381 4408 443
rect 4470 381 4504 443
rect 4566 381 4602 443
rect 4664 381 4698 443
rect 4752 353 4797 780
rect 3324 301 3330 353
rect 3382 350 3797 353
rect 4751 351 4797 353
rect 4599 350 4797 351
rect 3382 343 4797 350
rect 3382 308 3788 343
rect 3382 301 3388 308
rect 3786 287 3788 308
rect 3841 308 3980 343
rect 3841 287 3842 308
rect 3786 280 3842 287
rect 3978 287 3980 308
rect 4033 308 4172 343
rect 4033 287 4034 308
rect 3978 280 4034 287
rect 4170 287 4172 308
rect 4225 308 4364 343
rect 4225 287 4226 308
rect 4170 280 4226 287
rect 4362 287 4364 308
rect 4417 308 4556 343
rect 4417 287 4418 308
rect 4362 280 4418 287
rect 4554 287 4556 308
rect 4609 308 4797 343
rect 4609 287 4611 308
rect 4554 280 4611 287
rect 2468 210 2808 280
rect 1142 -560 1212 210
rect 2603 -281 2673 210
rect 2603 -560 2673 -418
rect 4064 -560 4134 210
rect 1142 -630 4134 -560
use ota_bias  ota_bias_0
timestamp 1668153059
transform 1 0 2638 0 1 -350
box -551 -280 551 280
use ota_half  ota_half_0
timestamp 1668153059
transform 1 0 53 0 1 613
box -53 -613 2585 525
use ota_half  ota_half_1
timestamp 1668153059
transform -1 0 5223 0 1 613
box -53 -613 2585 525
<< labels >>
rlabel metal2 0 849 70 919 0 vdd
port 1 n
rlabel metal2 1142 -630 1212 -560 0 vss
port 2 n
rlabel metal1 2365 -248 2911 -202 5 vbias
port 5 n
rlabel metal2 4752 524 4797 596 0 out
port 6 n
rlabel metal2 2603 -70 2673 0 0 net1
rlabel metal1 2168 132 2330 178 7 in_n
port 4 n
rlabel metal1 2946 132 3108 178 3 in_p
port 3 n
<< end >>
