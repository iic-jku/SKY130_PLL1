magic
tech sky130A
magscale 1 2
timestamp 1661273666
<< metal1 >>
rect 1711 1811 1763 1817
rect 1711 1753 1763 1759
rect 1540 1436 1582 1528
rect 1711 1342 1763 1348
rect 1711 1284 1763 1290
rect 1720 1164 1754 1284
rect 2548 854 2582 1852
rect 1711 -237 1763 -231
rect 1711 -295 1763 -289
rect 1540 -612 1582 -520
rect 1711 -706 1763 -700
rect 1711 -764 1763 -758
rect 1720 -884 1754 -764
rect 2548 -1194 2582 -196
rect 1720 -2712 1754 -2340
rect 2139 -3054 2181 -2568
rect 2548 -2904 2582 -2244
<< via1 >>
rect 1711 1759 1763 1811
rect 1711 1290 1763 1342
rect 1711 -289 1763 -237
rect 1711 -758 1763 -706
<< metal2 >>
rect 1498 3019 1540 3061
rect 2720 3019 2762 3061
rect 1705 1759 1711 1811
rect 1763 1759 1769 1811
rect 1720 1342 1754 1759
rect 1705 1290 1711 1342
rect 1763 1290 1769 1342
rect 1498 971 1540 1013
rect 2720 971 2762 1013
rect 1705 -289 1711 -237
rect 1763 -289 1769 -237
rect 1720 -706 1754 -289
rect 1705 -758 1711 -706
rect 1763 -758 1769 -706
rect 1498 -1077 1540 -1035
rect 2720 -1077 2762 -1035
rect 1801 -2664 1843 -2388
rect 2468 -2856 2510 -2292
rect 2468 -3478 2510 -3298
rect 1801 -3670 1843 -3490
use tgate_1  tgate_1_0
timestamp 1660934390
transform 1 0 1801 0 1 2480
box -261 -952 919 1138
use tgate_1  tgate_1_1
timestamp 1660934390
transform 1 0 1801 0 1 432
box -261 -952 919 1138
use tgate_1  tgate_1_2
timestamp 1660934390
transform 1 0 1801 0 1 -1616
box -261 -952 919 1138
use vc_1  vc_1_0
timestamp 1660924909
transform 0 -1 2107 1 0 -3575
box -53 -613 1049 525
<< labels >>
rlabel metal2 2720 -1077 2762 -1035 0 b0
rlabel metal2 2720 971 2762 1013 6 b1
rlabel metal2 2720 3019 2762 3061 0 b2
rlabel metal2 2468 -3478 2510 -3436 7 vss
rlabel metal2 1801 -3670 1843 -3628 7 vdd
rlabel metal2 1498 -1077 1540 -1035 1 ss
rlabel metal2 1498 971 1540 1013 0 tt
rlabel metal2 1498 3019 1540 3061 0 ff
<< end >>
