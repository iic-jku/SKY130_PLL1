magic
tech sky130A
magscale 1 2
timestamp 1659991419
<< error_s >>
rect -121 387 -63 393
rect 1127 387 1185 393
rect 1811 387 1869 393
rect 2867 387 2925 393
rect 3551 387 3609 393
rect 4415 387 4473 393
rect -121 353 -109 387
rect 1127 353 1139 387
rect 1811 353 1823 387
rect 2867 353 2879 387
rect 3551 353 3563 387
rect 4415 353 4427 387
rect -121 347 -63 353
rect 1127 347 1185 353
rect 1811 347 1869 353
rect 2867 347 2925 353
rect 3551 347 3609 353
rect 4415 347 4473 353
rect -121 -459 -63 -453
rect 1127 -459 1185 -453
rect 1811 -459 1869 -453
rect 2867 -459 2925 -453
rect -121 -493 -109 -459
rect 1127 -493 1139 -459
rect 1811 -493 1823 -459
rect 2867 -493 2879 -459
rect -121 -499 -63 -493
rect 1127 -499 1185 -493
rect 1811 -499 1869 -493
rect 2867 -499 2925 -493
rect 455 -1019 513 -1013
rect 1127 -1019 1185 -1013
rect 1811 -1019 1869 -1013
rect 2291 -1019 2349 -1013
rect 3551 -1019 3609 -1013
rect 4031 -1019 4089 -1013
rect 455 -1053 467 -1019
rect 1127 -1053 1139 -1019
rect 1811 -1053 1823 -1019
rect 2291 -1053 2303 -1019
rect 3551 -1053 3563 -1019
rect 4031 -1053 4043 -1019
rect 455 -1059 513 -1053
rect 1127 -1059 1185 -1053
rect 1811 -1059 1869 -1053
rect 2291 -1059 2349 -1053
rect 3551 -1059 3609 -1053
rect 4031 -1059 4089 -1053
rect 1811 -1329 1869 -1323
rect 2291 -1329 2349 -1323
rect 3551 -1329 3609 -1323
rect 4031 -1329 4089 -1323
rect 1811 -1363 1823 -1329
rect 2291 -1363 2303 -1329
rect 3551 -1363 3563 -1329
rect 4031 -1363 4043 -1329
rect 1811 -1369 1869 -1363
rect 2291 -1369 2349 -1363
rect 3551 -1369 3609 -1363
rect 4031 -1369 4089 -1363
<< locali >>
rect 627 -1548 659 -1514
rect 693 -1548 755 -1514
rect 789 -1548 831 -1514
<< viali >>
rect 659 -1548 693 -1514
rect 755 -1548 789 -1514
<< metal1 >>
rect 1371 119 1377 128
rect 1089 85 1377 119
rect 1371 76 1377 85
rect 1429 76 1435 128
rect 1481 76 1487 128
rect 1539 119 1545 128
rect 1539 85 1907 119
rect 1539 76 1545 85
rect 3232 76 3238 128
rect 3290 119 3296 128
rect 3290 85 3647 119
rect 3290 76 3296 85
rect -307 -225 -25 -191
rect 1089 -225 1907 -191
rect 1371 -769 1377 -760
rect 1089 -803 1377 -769
rect 1371 -812 1377 -803
rect 1429 -812 1435 -760
rect 1591 -769 1625 -225
rect 1591 -803 1907 -769
rect 2253 -803 3647 -769
rect 705 -1376 711 -1367
rect 664 -1410 711 -1376
rect 705 -1419 711 -1410
rect 763 -1419 769 -1367
rect 644 -1514 650 -1505
rect 702 -1514 708 -1505
rect 740 -1514 746 -1505
rect 798 -1514 804 -1505
rect 627 -1548 650 -1514
rect 702 -1548 746 -1514
rect 798 -1548 831 -1514
rect 644 -1557 650 -1548
rect 702 -1557 708 -1548
rect 740 -1557 746 -1548
rect 798 -1557 804 -1548
rect 1481 -1622 1487 -1570
rect 1539 -1579 1545 -1570
rect 1539 -1613 1907 -1579
rect 1539 -1622 1545 -1613
rect 3232 -1622 3238 -1570
rect 3290 -1579 3296 -1570
rect 3290 -1613 3647 -1579
rect 3290 -1622 3296 -1613
<< via1 >>
rect 1377 76 1429 128
rect 1487 76 1539 128
rect 3238 76 3290 128
rect 1377 -812 1429 -760
rect 711 -1419 763 -1367
rect 650 -1514 702 -1505
rect 746 -1514 798 -1505
rect 650 -1548 659 -1514
rect 659 -1548 693 -1514
rect 693 -1548 702 -1514
rect 746 -1548 755 -1514
rect 755 -1548 789 -1514
rect 789 -1548 798 -1514
rect 650 -1557 702 -1548
rect 746 -1557 798 -1548
rect 1487 -1622 1539 -1570
rect 3238 -1622 3290 -1570
<< metal2 >>
rect 502 -272 562 166
rect 1377 128 1429 134
rect 1377 70 1429 76
rect 1487 128 1539 134
rect 1487 70 1539 76
rect 1386 -38 1420 70
rect 1376 -47 1432 -38
rect 1376 -112 1432 -103
rect 502 -492 562 -483
rect 502 -561 562 -552
rect 510 -609 554 -561
rect 510 -653 842 -609
rect 798 -842 842 -653
rect 1386 -754 1420 -112
rect 1496 -345 1530 70
rect 2338 -272 2398 166
rect 3238 128 3290 134
rect 3238 70 3290 76
rect 3247 -345 3281 70
rect 3792 -47 3848 -38
rect 3990 -53 4034 166
rect 3848 -97 4034 -53
rect 3792 -112 3848 -103
rect 1485 -354 1541 -345
rect 1485 -419 1541 -410
rect 3236 -354 3292 -345
rect 3236 -419 3292 -410
rect 1377 -760 1429 -754
rect 1377 -818 1429 -812
rect 720 -1361 754 -1332
rect 711 -1367 763 -1361
rect 711 -1425 763 -1419
rect 143 -1446 203 -1437
rect 702 -1499 746 -1478
rect 143 -1515 203 -1506
rect 650 -1505 798 -1499
rect 151 -1572 195 -1515
rect 702 -1557 746 -1505
rect 650 -1563 798 -1557
rect 1496 -1564 1530 -419
rect 2058 -1401 2102 -981
rect 3247 -1564 3281 -419
rect 3798 -557 3842 -112
rect 3790 -566 3850 -557
rect 3790 -635 3850 -626
rect 3798 -1401 3842 -981
rect 1487 -1570 1539 -1564
rect 1487 -1628 1539 -1622
rect 3238 -1570 3290 -1564
rect 3238 -1628 3290 -1622
<< via2 >>
rect 1376 -103 1432 -47
rect 502 -552 562 -492
rect 3792 -103 3848 -47
rect 1485 -410 1541 -354
rect 3236 -410 3292 -354
rect 143 -1506 203 -1446
rect 3790 -626 3850 -566
<< metal3 >>
rect -307 246 -177 306
rect 1241 246 1755 306
rect 2981 246 3495 306
rect 4529 246 4659 306
rect 1371 -45 1437 -42
rect 3787 -45 3853 -42
rect 1371 -47 4659 -45
rect 1371 -103 1376 -47
rect 1432 -103 3792 -47
rect 3848 -103 4659 -47
rect 1371 -105 4659 -103
rect 1371 -108 1437 -105
rect 3787 -108 3853 -105
rect 1480 -352 1546 -349
rect 3231 -352 3297 -349
rect 1241 -354 1546 -352
rect 1241 -410 1485 -354
rect 1541 -410 1546 -354
rect 1241 -412 1546 -410
rect 2981 -354 3297 -352
rect 2981 -410 3236 -354
rect 3292 -410 3297 -354
rect 2981 -412 3297 -410
rect 502 -487 562 -414
rect 1480 -415 1546 -412
rect 2309 -414 2427 -412
rect 497 -492 567 -487
rect 497 -552 502 -492
rect 562 -552 567 -492
rect 497 -557 567 -552
rect 2338 -601 2398 -414
rect 3231 -415 3297 -412
rect 2050 -661 2398 -601
rect 3785 -566 3855 -561
rect 3785 -626 3790 -566
rect 3850 -626 3855 -566
rect 3785 -631 3855 -626
rect 2050 -839 2110 -661
rect 3790 -839 3850 -631
rect 1241 -981 1431 -921
rect 143 -1441 203 -1278
rect 138 -1446 208 -1441
rect 138 -1506 143 -1446
rect 203 -1506 208 -1446
rect 138 -1511 208 -1506
rect 1370 -1481 1430 -981
rect 1370 -1541 1755 -1481
rect 2405 -1541 3495 -1481
rect 4145 -1541 4275 -1481
use d_ff_n2  sky130_fd_pr__nfet_01v8_GVQ53W_0
timestamp 1659939748
transform 1 0 2080 0 1 -911
box -525 -280 455 280
use d_ff_n2  sky130_fd_pr__nfet_01v8_GVQ53W_1
timestamp 1659939748
transform -1 0 2080 0 -1 -1471
box -525 -280 455 280
use d_ff_n2  sky130_fd_pr__nfet_01v8_GVQ53W_2
timestamp 1659939748
transform 1 0 3820 0 1 -911
box -525 -280 455 280
use d_ff_n2  sky130_fd_pr__nfet_01v8_GVQ53W_3
timestamp 1659939748
transform -1 0 3820 0 -1 -1471
box -525 -280 455 280
use d_ff_n1  sky130_fd_pr__nfet_01v8_WWA63A_0
timestamp 1659940462
transform 1 0 820 0 1 -911
box -551 -280 621 280
use d_ff_p2  sky130_fd_pr__pfet_01v8_BD2UMN_0
timestamp 1659939748
transform 1 0 2368 0 1 236
box -813 -289 743 289
use d_ff_p2  sky130_fd_pr__pfet_01v8_BD2UMN_1
timestamp 1659939748
transform -1 0 2368 0 -1 -342
box -813 -289 743 289
use d_ff_p3  sky130_fd_pr__pfet_01v8_BDAGKN_0
timestamp 1659939748
transform 1 0 4012 0 1 236
box -647 -289 717 289
use d_ff_p1  sky130_fd_pr__pfet_01v8_BDS2ZN_0
timestamp 1659940462
transform 1 0 532 0 1 236
box -909 -289 839 289
use d_ff_p1  sky130_fd_pr__pfet_01v8_BDS2ZN_1
timestamp 1659940462
transform -1 0 532 0 -1 -342
box -909 -289 839 289
<< end >>
