magic
tech sky130A
magscale 1 2
timestamp 1668431035
<< nwell >>
rect 6655 -68 7423 498
rect 9402 476 10253 1042
rect 9402 -612 10258 -46
<< pwell >>
rect 9449 1146 9930 1282
rect 4974 602 5458 738
rect -85 21 4577 157
rect 9449 236 9930 372
rect 9449 58 9930 194
rect 4976 -308 5458 -172
rect 9449 -852 9930 -716
<< psubdiff >>
rect 9614 1250 9910 1256
rect 9614 1178 9641 1250
rect 9878 1178 9910 1250
rect 9614 1169 9910 1178
rect 4999 704 5289 711
rect 4999 641 5024 704
rect 5263 641 5289 704
rect 4999 634 5289 641
rect 9614 349 9910 358
rect 9614 277 9641 349
rect 9878 277 9910 349
rect 9614 271 9910 277
rect 9614 169 9910 175
rect 1045 99 1296 108
rect 1045 60 1073 99
rect 1271 60 1296 99
rect 9614 97 9641 169
rect 9878 97 9910 169
rect 9614 88 9910 97
rect 1045 54 1296 60
rect 4994 -203 5290 -194
rect 4994 -275 5021 -203
rect 5258 -275 5290 -203
rect 4994 -281 5290 -275
rect 9613 -749 9909 -740
rect 9613 -821 9640 -749
rect 9877 -821 9909 -749
rect 9613 -827 9909 -821
<< nsubdiff >>
rect 9971 825 10111 860
rect 9971 698 9981 825
rect 10099 698 10111 825
rect 9971 664 10111 698
rect 2311 475 2401 499
rect 2311 326 2322 475
rect 2389 326 2401 475
rect 2311 302 2401 326
rect 7246 282 7386 317
rect 7246 155 7256 282
rect 7374 155 7386 282
rect 7246 121 7386 155
rect 9971 -263 10111 -228
rect 9971 -390 9981 -263
rect 10099 -390 10111 -263
rect 9971 -424 10111 -390
<< psubdiffcont >>
rect 9641 1178 9878 1250
rect 5024 641 5263 704
rect 9641 277 9878 349
rect 1073 60 1271 99
rect 9641 97 9878 169
rect 5021 -275 5258 -203
rect 9640 -821 9877 -749
<< nsubdiffcont >>
rect 9981 698 10099 825
rect 2322 326 2389 475
rect 7256 155 7374 282
rect 9981 -390 10099 -263
<< poly >>
rect 1652 215 1747 249
rect 2775 222 2842 256
<< locali >>
rect 9595 1287 9934 1321
rect 9623 1250 9900 1287
rect 9623 1178 9641 1250
rect 9878 1178 9900 1250
rect 9623 1169 9900 1178
rect 9977 825 10104 841
rect 9977 780 9981 825
rect 5003 704 5280 776
rect 9904 737 9981 780
rect 5003 641 5024 704
rect 5263 641 5280 704
rect 9977 698 9981 737
rect 10099 698 10104 825
rect 9977 682 10104 698
rect 5003 634 5280 641
rect 2296 527 2436 561
rect 2296 475 2429 527
rect 2296 326 2322 475
rect 2389 326 2429 475
rect 9623 349 9900 358
rect 1011 313 1067 326
rect 1011 153 1023 313
rect 1057 153 1067 313
rect 2198 307 2254 320
rect 1264 249 2137 255
rect 1264 215 1271 249
rect 2128 215 2137 249
rect 1264 210 2137 215
rect 1011 145 1067 153
rect 2198 147 2210 307
rect 2244 147 2254 307
rect 2296 303 2429 326
rect 2296 302 2424 303
rect 7252 282 7379 298
rect 7252 237 7256 282
rect 7156 194 7256 237
rect 2198 139 2254 147
rect 7252 155 7256 194
rect 7374 155 7379 282
rect 9623 277 9641 349
rect 9878 277 9900 349
rect 9623 240 9900 277
rect 9595 206 9934 240
rect 7252 139 7379 155
rect 9623 169 9900 206
rect 1056 99 1287 105
rect 1056 60 1073 99
rect 1271 60 1287 99
rect 9623 97 9641 169
rect 9878 97 9900 169
rect 9623 88 9900 97
rect 1056 17 1287 60
rect 1059 -18 1285 17
rect 5003 -203 5280 -194
rect 5003 -275 5021 -203
rect 5258 -275 5280 -203
rect 5003 -346 5280 -275
rect 9977 -263 10104 -247
rect 9977 -308 9981 -263
rect 9904 -351 9981 -308
rect 9977 -390 9981 -351
rect 10099 -390 10104 -263
rect 9977 -406 10104 -390
rect 9622 -749 9899 -740
rect 9622 -821 9640 -749
rect 9877 -821 9899 -749
rect 9622 -858 9899 -821
rect 9594 -892 9933 -858
<< viali >>
rect 7823 1054 7988 1088
rect 8363 962 8397 996
rect 8535 962 8569 996
rect 8720 962 8773 996
rect 8917 962 8951 996
rect 9089 962 9123 996
rect 9261 962 9295 996
rect 5076 510 5241 544
rect 8362 522 8396 556
rect 8534 522 8568 556
rect 8719 522 8772 556
rect 8916 522 8950 556
rect 9088 522 9122 556
rect 9260 522 9294 556
rect 5616 418 5650 452
rect 5788 418 5822 452
rect 5973 418 6026 452
rect 6170 418 6204 452
rect 6342 418 6376 452
rect 6514 418 6548 452
rect 7823 429 7988 464
rect 9763 430 9841 465
rect 47 216 217 250
rect 307 153 341 313
rect 540 218 967 252
rect 1023 153 1057 313
rect 1271 215 2128 249
rect 2210 147 2244 307
rect 3075 307 3109 341
rect 3247 307 3281 341
rect 3432 307 3485 341
rect 3629 307 3663 341
rect 3801 307 3835 341
rect 3973 307 4007 341
rect 2536 209 2701 249
rect 4469 215 4544 249
rect 5615 -22 5649 12
rect 5787 -22 5821 12
rect 5972 -22 6025 12
rect 6169 -22 6203 12
rect 6341 -22 6375 12
rect 6513 -22 6547 12
rect 7823 -34 7988 0
rect 5076 -115 5241 -80
rect 7016 -114 7094 -79
rect 8363 -126 8397 -92
rect 8535 -126 8569 -92
rect 8720 -126 8773 -92
rect 8917 -126 8951 -92
rect 9089 -126 9123 -92
rect 9261 -126 9295 -92
rect 8362 -566 8396 -532
rect 8534 -566 8568 -532
rect 8719 -566 8772 -532
rect 8916 -566 8950 -532
rect 9088 -566 9122 -532
rect 9260 -566 9294 -532
rect 7823 -659 7988 -624
rect 9763 -658 9841 -623
<< metal1 >>
rect 5769 1617 6235 1623
rect 37 1421 503 1427
rect 37 721 503 955
rect 3999 1421 4465 1427
rect 3999 721 4465 955
rect 7722 1470 9929 1480
rect 7722 1450 9930 1470
rect 7722 1277 7744 1450
rect 9899 1277 9930 1450
rect 7722 1255 9930 1277
rect 5769 936 6235 1151
rect 7469 1088 8166 1215
rect -111 496 4644 721
rect 4975 711 7183 936
rect 4722 544 5419 671
rect 4722 446 4937 544
rect 5043 510 5076 544
rect 5241 510 5419 544
rect 5043 495 5419 510
rect 4034 383 4937 446
rect 3063 346 4937 383
rect 5604 452 6675 476
rect 5604 418 5616 452
rect 5650 418 5788 452
rect 5822 418 5973 452
rect 6026 418 6170 452
rect 6204 418 6342 452
rect 6376 418 6514 452
rect 6548 418 6675 452
rect 5604 413 6675 418
rect 7469 429 7684 1088
rect 7790 1054 7823 1088
rect 7988 1054 8166 1088
rect 7790 1039 8166 1054
rect 8351 996 9422 1020
rect 8351 962 8363 996
rect 8397 962 8535 996
rect 8569 962 8720 996
rect 8773 962 8917 996
rect 8951 962 9089 996
rect 9123 962 9261 996
rect 9295 962 9422 996
rect 8351 957 9422 962
rect 8351 920 10254 957
rect 9322 857 10254 920
rect 7722 788 7890 807
rect 7722 728 7737 788
rect 7722 711 7890 728
rect 10039 661 10254 857
rect 9321 598 10254 661
rect 8350 561 10254 598
rect 8350 556 9421 561
rect 8350 522 8362 556
rect 8396 522 8534 556
rect 8568 522 8719 556
rect 8772 522 8916 556
rect 8950 522 9088 556
rect 9122 522 9260 556
rect 9294 522 9421 556
rect 8350 498 9421 522
rect 7790 464 8165 476
rect 7790 429 7823 464
rect 7988 429 8165 464
rect 7469 413 8165 429
rect 5604 376 8165 413
rect 9507 465 9864 476
rect 9507 430 9763 465
rect 9841 430 9864 465
rect 9507 394 9864 430
rect 10039 449 10254 561
rect 3063 341 4134 346
rect -184 250 261 326
rect -184 216 47 250
rect 217 216 261 250
rect -184 145 261 216
rect 295 313 976 326
rect 295 153 307 313
rect 341 252 976 313
rect 341 218 540 252
rect 967 218 976 252
rect 341 153 976 218
rect 295 145 976 153
rect 1011 324 1236 326
rect 1011 313 2137 324
rect 1011 153 1023 313
rect 1057 249 2137 313
rect 1057 215 1271 249
rect 2128 215 2137 249
rect 1057 153 2137 215
rect 1011 145 2137 153
rect 2198 307 2886 320
rect 2198 147 2210 307
rect 2244 249 2886 307
rect 3063 307 3075 341
rect 3109 307 3247 341
rect 3281 307 3432 341
rect 3485 307 3629 341
rect 3663 307 3801 341
rect 3835 307 3973 341
rect 4007 307 4134 341
rect 3063 283 4134 307
rect 2244 209 2536 249
rect 2701 209 2886 249
rect 2244 147 2886 209
rect 4222 249 4578 262
rect 4222 215 4469 249
rect 4544 215 4578 249
rect 4222 179 4578 215
rect 2198 139 2886 147
rect -115 -177 4644 48
rect 4722 -115 4937 346
rect 6575 313 8165 376
rect 7469 292 8165 313
rect 4975 244 5143 263
rect 4975 184 4990 244
rect 4975 167 5143 184
rect 7469 127 7684 292
rect 7722 244 7890 263
rect 7722 184 7737 244
rect 7722 167 7890 184
rect 7469 117 8166 127
rect 6574 54 8166 117
rect 5603 17 8166 54
rect 5603 12 6674 17
rect 5603 -22 5615 12
rect 5649 -22 5787 12
rect 5821 -22 5972 12
rect 6025 -22 6169 12
rect 6203 -22 6341 12
rect 6375 -22 6513 12
rect 6547 -22 6674 12
rect 5603 -46 6674 -22
rect 7469 0 8166 17
rect 5043 -80 5418 -68
rect 5043 -115 5076 -80
rect 5241 -115 5418 -80
rect 100 -329 566 -177
rect 100 -801 566 -795
rect 4000 -329 4466 -177
rect 4722 -252 5418 -115
rect 6760 -79 7117 -68
rect 6760 -114 7016 -79
rect 7094 -114 7117 -79
rect 6760 -150 7117 -114
rect 4975 -341 5787 -281
rect 6253 -341 7183 -281
rect 4975 -506 7183 -341
rect 4000 -801 4466 -795
rect 5787 -711 6253 -506
rect 7469 -659 7684 0
rect 7790 -34 7823 0
rect 7988 -34 8166 0
rect 7790 -49 8166 -34
rect 10039 -17 10797 449
rect 8351 -92 9422 -68
rect 8351 -126 8363 -92
rect 8397 -126 8535 -92
rect 8569 -126 8720 -92
rect 8773 -126 8917 -92
rect 8951 -126 9089 -92
rect 9123 -126 9261 -92
rect 9295 -126 9422 -92
rect 8351 -131 9422 -126
rect 10039 -131 10254 -17
rect 8351 -168 10254 -131
rect 9322 -231 10254 -168
rect 7722 -300 7890 -281
rect 7722 -360 7737 -300
rect 7722 -377 7890 -360
rect 10039 -427 10254 -231
rect 9321 -490 10254 -427
rect 8350 -527 10254 -490
rect 8350 -532 9421 -527
rect 8350 -566 8362 -532
rect 8396 -566 8534 -532
rect 8568 -566 8719 -532
rect 8772 -566 8916 -532
rect 8950 -566 9088 -532
rect 9122 -566 9260 -532
rect 9294 -566 9421 -532
rect 8350 -590 9421 -566
rect 7790 -624 8165 -612
rect 7790 -659 7823 -624
rect 7988 -659 8165 -624
rect 7469 -796 8165 -659
rect 9507 -623 9864 -612
rect 9507 -658 9763 -623
rect 9841 -658 9864 -623
rect 9507 -694 9864 -658
rect 7722 -846 9930 -825
rect 7722 -1019 7750 -846
rect 9905 -1019 9930 -846
rect 7722 -1050 9930 -1019
rect 5787 -1183 6253 -1177
<< via1 >>
rect 37 955 503 1421
rect 3999 955 4465 1421
rect 5769 1151 6235 1617
rect 7744 1277 9899 1450
rect 7737 728 9918 788
rect 4990 184 7171 244
rect 7737 184 9918 244
rect 100 -795 566 -329
rect 4000 -795 4466 -329
rect 5787 -1177 6253 -711
rect 7737 -360 9918 -300
rect 7750 -1019 9905 -846
<< metal2 >>
rect 7220 1982 7686 1991
rect 5769 1617 6235 1626
rect 37 1421 503 1430
rect 3999 1421 4465 1430
rect 31 955 37 1421
rect 503 955 509 1421
rect 3993 955 3999 1421
rect 4465 955 4471 1421
rect 5763 1151 5769 1617
rect 6235 1151 6241 1617
rect 5769 1142 6235 1151
rect 37 946 503 955
rect 3999 946 4465 955
rect 7220 807 7686 1516
rect 9992 1977 10458 1986
rect 9992 1480 10458 1511
rect 7722 1450 10458 1480
rect 7722 1277 7744 1450
rect 9899 1277 10458 1450
rect 7722 1255 10458 1277
rect 7220 788 9930 807
rect 7220 728 7737 788
rect 9918 728 9930 788
rect 7220 711 9930 728
rect 7220 263 7686 711
rect 9992 303 10458 1255
rect 9584 263 10458 303
rect 4975 244 7686 263
rect 4975 184 4990 244
rect 7171 184 7686 244
rect 4975 167 7686 184
rect 7722 244 10458 263
rect 7722 184 7737 244
rect 9918 184 10458 244
rect 7722 167 10458 184
rect 7220 -281 7686 167
rect 9584 128 10458 167
rect 7220 -300 9930 -281
rect 100 -329 566 -320
rect 4000 -329 4466 -320
rect 94 -795 100 -329
rect 566 -795 572 -329
rect 3994 -795 4000 -329
rect 4466 -795 4472 -329
rect 7220 -360 7737 -300
rect 9918 -360 9930 -300
rect 7220 -377 9930 -360
rect 5787 -711 6253 -702
rect 100 -804 566 -795
rect 4000 -804 4466 -795
rect 5781 -1177 5787 -711
rect 6253 -1177 6259 -711
rect 7220 -1109 7686 -377
rect 9992 -825 10458 128
rect 7722 -846 10458 -825
rect 7722 -1019 7750 -846
rect 9905 -1019 10458 -846
rect 7722 -1050 10458 -1019
rect 5787 -1186 6253 -1177
rect 9992 -1055 10458 -1050
rect 9992 -1530 10458 -1521
rect 7220 -1584 7686 -1575
<< via2 >>
rect 37 955 503 1421
rect 3999 955 4465 1421
rect 5769 1151 6235 1617
rect 7220 1516 7686 1982
rect 9992 1511 10458 1977
rect 100 -795 566 -329
rect 4000 -795 4466 -329
rect 5787 -1177 6253 -711
rect 7220 -1575 7686 -1109
rect 9992 -1521 10458 -1055
<< metal3 >>
rect 7215 1987 7691 1993
rect 5764 1622 6240 1628
rect 32 1426 508 1432
rect 32 955 37 960
rect 503 955 508 960
rect 32 950 508 955
rect 3994 1426 4470 1432
rect 7215 1516 7220 1521
rect 7686 1516 7691 1521
rect 7215 1511 7691 1516
rect 9987 1982 10463 1988
rect 9987 1511 9992 1516
rect 10458 1511 10463 1516
rect 9987 1506 10463 1511
rect 5764 1151 5769 1156
rect 6235 1151 6240 1156
rect 5764 1146 6240 1151
rect 3994 955 3999 960
rect 4465 955 4470 960
rect 3994 950 4470 955
rect 95 -329 571 -324
rect 95 -334 100 -329
rect 566 -334 571 -329
rect 95 -806 571 -800
rect 3995 -329 4471 -324
rect 3995 -334 4000 -329
rect 4466 -334 4471 -329
rect 3995 -806 4471 -800
rect 5782 -711 6258 -706
rect 5782 -716 5787 -711
rect 6253 -716 6258 -711
rect 9987 -1055 10463 -1050
rect 9987 -1060 9992 -1055
rect 10458 -1060 10463 -1055
rect 5782 -1188 6258 -1182
rect 7215 -1109 7691 -1104
rect 7215 -1114 7220 -1109
rect 7686 -1114 7691 -1109
rect 9987 -1532 10463 -1526
rect 7215 -1586 7691 -1580
<< via3 >>
rect 7215 1982 7691 1987
rect 5764 1617 6240 1622
rect 32 1421 508 1426
rect 32 960 37 1421
rect 37 960 503 1421
rect 503 960 508 1421
rect 3994 1421 4470 1426
rect 3994 960 3999 1421
rect 3999 960 4465 1421
rect 4465 960 4470 1421
rect 5764 1156 5769 1617
rect 5769 1156 6235 1617
rect 6235 1156 6240 1617
rect 7215 1521 7220 1982
rect 7220 1521 7686 1982
rect 7686 1521 7691 1982
rect 9987 1977 10463 1982
rect 9987 1516 9992 1977
rect 9992 1516 10458 1977
rect 10458 1516 10463 1977
rect 95 -795 100 -334
rect 100 -795 566 -334
rect 566 -795 571 -334
rect 95 -800 571 -795
rect 3995 -795 4000 -334
rect 4000 -795 4466 -334
rect 4466 -795 4471 -334
rect 3995 -800 4471 -795
rect 5782 -1177 5787 -716
rect 5787 -1177 6253 -716
rect 6253 -1177 6258 -716
rect 5782 -1182 6258 -1177
rect 7215 -1575 7220 -1114
rect 7220 -1575 7686 -1114
rect 7686 -1575 7691 -1114
rect 9987 -1521 9992 -1060
rect 9992 -1521 10458 -1060
rect 10458 -1521 10463 -1060
rect 9987 -1526 10463 -1521
rect 7215 -1580 7691 -1575
<< metal4 >>
rect -276 2070 10919 2293
rect -276 1987 9879 2070
rect -276 1723 7215 1987
rect -276 1426 5665 1723
rect -276 960 32 1426
rect 508 960 3994 1426
rect 4470 1062 5665 1426
rect 5763 1156 5764 1157
rect 6240 1156 6241 1157
rect 5763 1155 6241 1156
rect 6362 1521 7215 1723
rect 7691 1521 9879 1987
rect 6362 1409 9879 1521
rect 9986 1516 9987 1517
rect 10463 1516 10464 1517
rect 9986 1515 10464 1516
rect 10576 1409 10919 2070
rect 6362 1062 10919 1409
rect 4470 960 10919 1062
rect -276 -230 10919 960
rect -276 -891 -16 -230
rect 681 -238 10919 -230
rect 94 -334 572 -333
rect 94 -335 95 -334
rect 571 -335 572 -334
rect 681 -891 3886 -238
rect 3994 -334 4472 -333
rect 3994 -335 3995 -334
rect 4471 -335 4472 -334
rect 4583 -613 10919 -238
rect -276 -899 3886 -891
rect 4583 -899 5676 -613
rect -276 -1274 5676 -899
rect 5781 -716 6259 -715
rect 5781 -717 5782 -716
rect 6258 -717 6259 -716
rect 6373 -943 10919 -613
rect 6373 -1114 9876 -943
rect 6373 -1274 7215 -1114
rect -276 -1580 7215 -1274
rect 7691 -1580 9876 -1114
rect 9986 -1060 10464 -1059
rect 9986 -1061 9987 -1060
rect 10463 -1061 10464 -1060
rect -276 -1604 9876 -1580
rect 10573 -1604 10919 -943
rect -276 -1892 10919 -1604
<< via4 >>
rect 5763 1622 6241 1623
rect 5763 1157 5764 1622
rect 5764 1157 6240 1622
rect 6240 1157 6241 1622
rect 9986 1982 10464 1983
rect 9986 1517 9987 1982
rect 9987 1517 10463 1982
rect 10463 1517 10464 1982
rect 94 -800 95 -335
rect 95 -800 571 -335
rect 571 -800 572 -335
rect 94 -801 572 -800
rect 3994 -800 3995 -335
rect 3995 -800 4471 -335
rect 4471 -800 4472 -335
rect 3994 -801 4472 -800
rect 5781 -1182 5782 -717
rect 5782 -1182 6258 -717
rect 6258 -1182 6259 -717
rect 5781 -1183 6259 -1182
rect 9986 -1526 9987 -1061
rect 9987 -1526 10463 -1061
rect 10463 -1526 10464 -1061
rect 9986 -1527 10464 -1526
<< metal5 >>
rect -276 1983 10919 2293
rect -276 1623 9986 1983
rect -276 1157 5763 1623
rect 6241 1517 9986 1623
rect 10464 1517 10919 1983
rect 6241 1157 10919 1517
rect -276 -335 10919 1157
rect -276 -801 94 -335
rect 572 -801 3994 -335
rect 4472 -717 10919 -335
rect 4472 -801 5781 -717
rect -276 -1183 5781 -801
rect 6259 -1061 10919 -717
rect 6259 -1183 9986 -1061
rect -276 -1527 9986 -1183
rect 10464 -1527 10919 -1061
rect -276 -1892 10919 -1527
use sky130_fd_sc_hd__clkinv_2  sky130_fd_sc_hd__clkinv_2_0 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 0 0 1 0
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_4  sky130_fd_sc_hd__clkinv_4_0 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 444 0 1 0
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_8  sky130_fd_sc_hd__clkinv_8_0 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1164 0 1 0
box -38 -48 1234 592
use sky130_fd_sc_hd__clkinv_16  sky130_fd_sc_hd__clkinv_16_0 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 2436 0 1 0
box -38 -48 2246 592
use sky130_fd_sc_hd__clkinv_16  sky130_fd_sc_hd__clkinv_16_1
timestamp 1666464484
transform 1 0 7722 0 -1 215
box -38 -48 2246 592
use sky130_fd_sc_hd__clkinv_16  sky130_fd_sc_hd__clkinv_16_2
timestamp 1666464484
transform 1 0 4975 0 -1 759
box -38 -48 2246 592
use sky130_fd_sc_hd__clkinv_16  sky130_fd_sc_hd__clkinv_16_3
timestamp 1666464484
transform 1 0 4975 0 1 -329
box -38 -48 2246 592
use sky130_fd_sc_hd__clkinv_16  sky130_fd_sc_hd__clkinv_16_4
timestamp 1666464484
transform 1 0 7722 0 1 -873
box -38 -48 2246 592
use sky130_fd_sc_hd__clkinv_16  sky130_fd_sc_hd__clkinv_16_5
timestamp 1666464484
transform 1 0 7722 0 1 215
box -38 -48 2246 592
use sky130_fd_sc_hd__clkinv_16  sky130_fd_sc_hd__clkinv_16_6
timestamp 1666464484
transform 1 0 7722 0 -1 1303
box -38 -48 2246 592
<< labels >>
rlabel metal1 -184 145 -3 326 3 in
port 3 n
rlabel metal1 10039 106 10254 322 0 out
port 4 n
rlabel metal1 -110 496 -14 592 7 vdd
rlabel metal1 -115 -48 -19 48 0 vss
rlabel metal2 7220 -1430 7686 -964 0 vdd
port 1 n
rlabel metal2 9992 -1512 10458 -1046 0 vss
port 2 n
rlabel metal1 5769 904 6235 1370 0 vss
rlabel metal1 5787 -929 6253 -463 0 vss
rlabel metal1 4000 -544 4466 -78 7 vss
rlabel metal1 100 -544 566 -78 7 vss
rlabel metal1 3999 629 4465 1095 7 vdd
rlabel metal1 37 629 503 1095 7 vdd
<< end >>
