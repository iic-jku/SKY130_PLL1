magic
tech sky130A
timestamp 1654412581
<< nwell >>
rect -251 -144 251 144
<< pmos >>
rect -151 -35 -136 35
rect -103 -35 -88 35
rect -55 -35 -40 35
rect -7 -35 7 35
rect 40 -35 55 35
rect 88 -35 103 35
rect 136 -35 151 35
<< pdiff >>
rect -182 29 -151 35
rect -182 -29 -176 29
rect -159 -29 -151 29
rect -182 -35 -151 -29
rect -136 29 -103 35
rect -136 -29 -128 29
rect -111 -29 -103 29
rect -136 -35 -103 -29
rect -88 29 -55 35
rect -88 -29 -80 29
rect -63 -29 -55 29
rect -88 -35 -55 -29
rect -40 29 -7 35
rect -40 -29 -32 29
rect -15 -29 -7 29
rect -40 -35 -7 -29
rect 7 29 40 35
rect 7 -29 15 29
rect 32 -29 40 29
rect 7 -35 40 -29
rect 55 29 88 35
rect 55 -29 63 29
rect 80 -29 88 29
rect 55 -35 88 -29
rect 103 29 136 35
rect 103 -29 111 29
rect 128 -29 136 29
rect 103 -35 136 -29
rect 151 29 182 35
rect 151 -29 159 29
rect 176 -29 182 29
rect 151 -35 182 -29
<< pdiffc >>
rect -176 -29 -159 29
rect -128 -29 -111 29
rect -80 -29 -63 29
rect -32 -29 -15 29
rect 15 -29 32 29
rect 63 -29 80 29
rect 111 -29 128 29
rect 159 -29 176 29
<< nsubdiff >>
rect -233 109 -185 126
rect 185 109 233 126
rect -233 78 -216 109
rect 216 78 233 109
rect -233 -109 -216 -78
rect 216 -109 233 -78
rect -233 -126 -185 -109
rect 185 -126 233 -109
<< nsubdiffcont >>
rect -185 109 185 126
rect -233 -78 -216 78
rect 216 -78 233 78
rect -185 -126 185 -109
<< poly >>
rect -112 75 16 83
rect -112 58 -104 75
rect -87 58 -56 75
rect -39 58 -8 75
rect 8 58 16 75
rect -112 50 16 58
rect 79 75 112 83
rect 79 58 87 75
rect 104 58 112 75
rect 79 50 112 58
rect -151 35 -136 48
rect -103 35 -88 50
rect -55 35 -40 50
rect -7 35 7 50
rect 40 35 55 48
rect 88 35 103 50
rect 136 35 151 48
rect -151 -50 -136 -35
rect -103 -48 -88 -35
rect -55 -48 -40 -35
rect -7 -48 7 -35
rect 40 -50 55 -35
rect 88 -48 103 -35
rect 136 -50 151 -35
rect -160 -58 -127 -50
rect -160 -75 -152 -58
rect -135 -75 -127 -58
rect -160 -83 -127 -75
rect 31 -58 64 -50
rect 31 -75 39 -58
rect 56 -75 64 -58
rect 31 -83 64 -75
rect 127 -58 160 -50
rect 127 -75 135 -58
rect 152 -75 160 -58
rect 127 -83 160 -75
<< polycont >>
rect -104 58 -87 75
rect -56 58 -39 75
rect -8 58 8 75
rect 87 58 104 75
rect -152 -75 -135 -58
rect 39 -75 56 -58
rect 135 -75 152 -58
<< locali >>
rect -233 109 -185 126
rect 185 109 233 126
rect -233 78 -216 109
rect 216 78 233 109
rect -112 58 -104 75
rect -87 58 -56 75
rect -39 58 -8 75
rect 8 58 16 75
rect 79 58 87 75
rect 104 58 112 75
rect -176 29 -159 37
rect -176 -37 -159 -29
rect -128 29 -111 37
rect -128 -37 -111 -29
rect -80 29 -63 37
rect -80 -37 -63 -29
rect -32 29 -15 37
rect -32 -37 -15 -29
rect 15 29 32 37
rect 15 -37 32 -29
rect 63 29 80 37
rect 63 -37 80 -29
rect 111 29 128 37
rect 111 -37 128 -29
rect 159 29 176 37
rect 159 -37 176 -29
rect -160 -75 -152 -58
rect -135 -75 -127 -58
rect 31 -75 39 -58
rect 56 -75 64 -58
rect 127 -75 135 -58
rect 152 -75 160 -58
rect -233 -109 -216 -78
rect 216 -109 233 -78
rect -233 -126 -185 -109
rect 185 -126 233 -109
<< viali >>
rect -104 58 -87 75
rect -56 58 -39 75
rect -8 58 8 75
rect 87 58 104 75
rect -176 -29 -159 29
rect -128 -29 -111 29
rect -80 -29 -63 29
rect -32 -29 -15 29
rect 15 -29 32 29
rect 63 -29 80 29
rect 111 -29 128 29
rect 159 -29 176 29
rect -152 -75 -135 -58
rect 39 -75 56 -58
rect 135 -75 152 -58
<< metal1 >>
rect -110 75 -81 78
rect -62 75 -33 78
rect -14 75 14 78
rect -251 58 -104 75
rect -87 58 -56 75
rect -39 58 -8 75
rect 8 58 14 75
rect -110 55 -81 58
rect -62 55 -33 58
rect -14 55 14 58
rect 81 75 110 78
rect 81 58 87 75
rect 104 58 128 75
rect 81 55 128 58
rect 111 35 128 55
rect -179 29 -156 35
rect -179 -29 -176 29
rect -159 -29 -156 29
rect -136 31 -103 35
rect -136 4 -133 31
rect -107 4 -103 31
rect -136 0 -128 4
rect -179 -35 -156 -29
rect -131 -29 -128 0
rect -111 0 -103 4
rect -83 29 -60 35
rect -83 0 -80 29
rect -111 -29 -108 0
rect -131 -35 -108 -29
rect -88 -5 -80 0
rect -63 0 -60 29
rect -40 31 -7 35
rect -40 4 -37 31
rect -11 4 -7 31
rect -40 0 -32 4
rect -63 -5 -55 0
rect -88 -32 -85 -5
rect -59 -32 -55 -5
rect -88 -35 -55 -32
rect -35 -29 -32 0
rect -15 0 -7 4
rect 12 29 35 35
rect 12 0 15 29
rect -15 -29 -12 0
rect -35 -35 -12 -29
rect 7 -5 15 0
rect 32 0 35 29
rect 55 31 88 35
rect 55 4 59 31
rect 85 4 88 31
rect 55 0 63 4
rect 32 -5 40 0
rect 7 -32 11 -5
rect 37 -32 40 -5
rect 7 -35 40 -32
rect 60 -29 63 0
rect 80 0 88 4
rect 108 29 131 35
rect 108 0 111 29
rect 80 -29 83 0
rect 60 -35 83 -29
rect 103 -5 111 0
rect 128 0 131 29
rect 156 29 179 35
rect 128 -5 136 0
rect 103 -32 107 -5
rect 133 -32 136 -5
rect 103 -35 136 -32
rect 156 -29 159 29
rect 176 -29 179 29
rect 156 -35 179 -29
rect 31 -54 64 -52
rect -158 -58 -129 -55
rect -158 -75 -152 -58
rect -135 -75 -43 -58
rect -158 -78 -129 -75
rect -61 -144 -43 -75
rect 31 -80 35 -54
rect 61 -80 64 -54
rect 129 -58 158 -55
rect 127 -75 135 -58
rect 152 -75 158 -58
rect 129 -78 158 -75
rect 31 -82 64 -80
rect 135 -144 152 -78
<< via1 >>
rect -133 29 -107 31
rect -133 4 -128 29
rect -128 4 -111 29
rect -111 4 -107 29
rect -37 29 -11 31
rect -37 4 -32 29
rect -32 4 -15 29
rect -15 4 -11 29
rect -85 -29 -80 -5
rect -80 -29 -63 -5
rect -63 -29 -59 -5
rect -85 -32 -59 -29
rect 59 29 85 31
rect 59 4 63 29
rect 63 4 80 29
rect 80 4 85 29
rect 11 -29 15 -5
rect 15 -29 32 -5
rect 32 -29 37 -5
rect 11 -32 37 -29
rect 107 -29 111 -5
rect 111 -29 128 -5
rect 128 -29 133 -5
rect 107 -32 133 -29
rect 35 -58 61 -54
rect 35 -75 39 -58
rect 39 -75 56 -58
rect 56 -75 61 -58
rect 35 -80 61 -75
<< metal2 >>
rect -138 32 -101 36
rect -138 3 -134 32
rect -106 3 -101 32
rect -138 -1 -101 3
rect -42 32 -5 36
rect -42 3 -38 32
rect -10 3 -5 32
rect -87 -5 -56 0
rect -42 -1 -5 3
rect 53 32 90 36
rect 53 3 58 32
rect 86 3 90 32
rect -87 -15 -85 -5
rect -251 -32 -85 -15
rect -59 -15 -56 -5
rect 9 -5 39 0
rect 53 -1 90 3
rect 9 -15 11 -5
rect -59 -32 11 -15
rect 37 -15 39 -5
rect 105 -5 135 0
rect 105 -15 107 -5
rect 37 -32 107 -15
rect 133 -32 135 -5
rect -251 -35 135 -32
rect 31 -54 64 -52
rect 31 -80 35 -54
rect 61 -80 64 -54
rect 31 -82 64 -80
rect 39 -144 56 -82
<< via2 >>
rect -134 31 -106 32
rect -134 4 -133 31
rect -133 4 -107 31
rect -107 4 -106 31
rect -134 3 -106 4
rect -38 31 -10 32
rect -38 4 -37 31
rect -37 4 -11 31
rect -11 4 -10 31
rect -38 3 -10 4
rect 58 31 86 32
rect 58 4 59 31
rect 59 4 85 31
rect 85 4 86 31
rect 58 3 86 4
<< metal3 >>
rect -91 37 -38 38
rect -251 32 251 37
rect -251 7 -134 32
rect -138 3 -134 7
rect -106 7 -38 32
rect -106 3 -101 7
rect -138 -1 -101 3
rect -42 3 -38 7
rect -10 7 58 32
rect -10 3 -5 7
rect -42 -1 -5 3
rect 53 3 58 7
rect 86 7 251 32
rect 86 3 90 7
rect 53 -1 90 3
<< properties >>
string FIXED_BBOX -225 -118 225 118
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.7 l 0.15 m 1 nf 7 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
