magic
tech sky130A
magscale 1 2
timestamp 1668109056
<< metal3 >>
rect -3186 66750 -1463 67041
rect 3185 66750 4908 67041
rect 9556 66750 11279 67041
rect 15927 66750 17650 67041
rect 22298 66750 24021 67041
rect -3186 62393 2894 66750
rect 3185 62393 9265 66750
rect 9556 62393 15636 66750
rect 15927 62393 22007 66750
rect 22298 62393 28378 66750
rect -3186 60670 28378 62393
rect -3186 60379 -1463 60670
rect 3185 60379 4908 60670
rect 9556 60379 11279 60670
rect 15927 60379 17650 60670
rect 22298 60379 24021 60670
rect -3186 56022 2894 60379
rect 3185 56022 9265 60379
rect 9556 56022 15636 60379
rect 15927 56022 22007 60379
rect 22298 56022 28378 60379
rect -3186 54299 28378 56022
rect -3186 54008 -1463 54299
rect 3185 54008 4908 54299
rect 9556 54008 11279 54299
rect 15927 54008 17650 54299
rect 22298 54008 24021 54299
rect -3186 49651 2894 54008
rect 3185 49651 9265 54008
rect 9556 49651 15636 54008
rect 15927 49651 22007 54008
rect 22298 49651 28378 54008
rect -3186 47928 28378 49651
rect -3186 47637 -1463 47928
rect 3185 47637 4908 47928
rect 9556 47637 11279 47928
rect 15927 47637 17650 47928
rect 22298 47637 24021 47928
rect -3186 43280 2894 47637
rect 3185 43280 9265 47637
rect 9556 43280 15636 47637
rect 15927 43280 22007 47637
rect 22298 43280 28378 47637
rect -3186 41557 28378 43280
rect -3186 41266 -1463 41557
rect 3185 41266 4908 41557
rect 9556 41266 11279 41557
rect 15927 41266 17650 41557
rect 22298 41266 24021 41557
rect -3186 36909 2894 41266
rect 3185 36909 9265 41266
rect 9556 36909 15636 41266
rect 15927 36909 22007 41266
rect 22298 36909 28378 41266
rect -3186 35186 28378 36909
rect -3186 34895 -1463 35186
rect 3185 34895 4908 35186
rect 9556 34895 11279 35186
rect 15927 34895 17650 35186
rect 22298 34895 24021 35186
rect -3186 30538 2894 34895
rect 3185 30538 9265 34895
rect 9556 30538 15636 34895
rect 15927 30538 22007 34895
rect 22298 30538 28378 34895
rect -3186 28815 28378 30538
rect -3186 28524 -1463 28815
rect 3185 28524 4908 28815
rect 9556 28524 11279 28815
rect 15927 28524 17650 28815
rect 22298 28524 24021 28815
rect -3186 24167 2894 28524
rect 3185 24167 9265 28524
rect 9556 24167 15636 28524
rect 15927 24167 22007 28524
rect 22298 24167 28378 28524
rect -3186 22444 28378 24167
rect -3186 22153 -1463 22444
rect 3185 22153 4908 22444
rect 9556 22153 11279 22444
rect 15927 22153 17650 22444
rect 22298 22153 24021 22444
rect -3186 17796 2894 22153
rect 3185 17796 9265 22153
rect 9556 17796 15636 22153
rect 15927 17796 22007 22153
rect 22298 17796 28378 22153
rect -3186 16073 28378 17796
rect -3186 15782 -1463 16073
rect 3185 15782 4908 16073
rect 9556 15782 11279 16073
rect 15927 15782 17650 16073
rect 22298 15782 24021 16073
rect -3186 11425 2894 15782
rect 3185 11425 9265 15782
rect 9556 11425 15636 15782
rect 15927 11425 22007 15782
rect 22298 11425 28378 15782
rect -3186 9702 28378 11425
rect -3186 9411 -1463 9702
rect 3185 9411 4908 9702
rect 9556 9411 11279 9702
rect 15927 9411 17650 9702
rect 22298 9411 24021 9702
rect -3186 5054 2894 9411
rect 3185 5054 9265 9411
rect 9556 5054 15636 9411
rect 15927 5054 22007 9411
rect 22298 5054 28378 9411
rect -3186 3331 28378 5054
rect -3186 3040 -1463 3331
rect 3185 3040 4908 3331
rect 9556 3040 11279 3331
rect 15927 3040 17650 3331
rect 22298 3040 24021 3331
rect -3186 -1317 2894 3040
rect 3185 -1317 9265 3040
rect 9556 -1317 15636 3040
rect 15927 -1317 22007 3040
rect 22298 -1317 28378 3040
rect -3186 -3040 28378 -1317
<< mimcap >>
rect -3146 66670 2854 66710
rect -3146 60750 -3106 66670
rect 2814 60750 2854 66670
rect -3146 60710 2854 60750
rect 3225 66670 9225 66710
rect 3225 60750 3265 66670
rect 9185 60750 9225 66670
rect 3225 60710 9225 60750
rect 9596 66670 15596 66710
rect 9596 60750 9636 66670
rect 15556 60750 15596 66670
rect 9596 60710 15596 60750
rect 15967 66670 21967 66710
rect 15967 60750 16007 66670
rect 21927 60750 21967 66670
rect 15967 60710 21967 60750
rect 22338 66670 28338 66710
rect 22338 60750 22378 66670
rect 28298 60750 28338 66670
rect 22338 60710 28338 60750
rect -3146 60299 2854 60339
rect -3146 54379 -3106 60299
rect 2814 54379 2854 60299
rect -3146 54339 2854 54379
rect 3225 60299 9225 60339
rect 3225 54379 3265 60299
rect 9185 54379 9225 60299
rect 3225 54339 9225 54379
rect 9596 60299 15596 60339
rect 9596 54379 9636 60299
rect 15556 54379 15596 60299
rect 9596 54339 15596 54379
rect 15967 60299 21967 60339
rect 15967 54379 16007 60299
rect 21927 54379 21967 60299
rect 15967 54339 21967 54379
rect 22338 60299 28338 60339
rect 22338 54379 22378 60299
rect 28298 54379 28338 60299
rect 22338 54339 28338 54379
rect -3146 53928 2854 53968
rect -3146 48008 -3106 53928
rect 2814 48008 2854 53928
rect -3146 47968 2854 48008
rect 3225 53928 9225 53968
rect 3225 48008 3265 53928
rect 9185 48008 9225 53928
rect 3225 47968 9225 48008
rect 9596 53928 15596 53968
rect 9596 48008 9636 53928
rect 15556 48008 15596 53928
rect 9596 47968 15596 48008
rect 15967 53928 21967 53968
rect 15967 48008 16007 53928
rect 21927 48008 21967 53928
rect 15967 47968 21967 48008
rect 22338 53928 28338 53968
rect 22338 48008 22378 53928
rect 28298 48008 28338 53928
rect 22338 47968 28338 48008
rect -3146 47557 2854 47597
rect -3146 41637 -3106 47557
rect 2814 41637 2854 47557
rect -3146 41597 2854 41637
rect 3225 47557 9225 47597
rect 3225 41637 3265 47557
rect 9185 41637 9225 47557
rect 3225 41597 9225 41637
rect 9596 47557 15596 47597
rect 9596 41637 9636 47557
rect 15556 41637 15596 47557
rect 9596 41597 15596 41637
rect 15967 47557 21967 47597
rect 15967 41637 16007 47557
rect 21927 41637 21967 47557
rect 15967 41597 21967 41637
rect 22338 47557 28338 47597
rect 22338 41637 22378 47557
rect 28298 41637 28338 47557
rect 22338 41597 28338 41637
rect -3146 41186 2854 41226
rect -3146 35266 -3106 41186
rect 2814 35266 2854 41186
rect -3146 35226 2854 35266
rect 3225 41186 9225 41226
rect 3225 35266 3265 41186
rect 9185 35266 9225 41186
rect 3225 35226 9225 35266
rect 9596 41186 15596 41226
rect 9596 35266 9636 41186
rect 15556 35266 15596 41186
rect 9596 35226 15596 35266
rect 15967 41186 21967 41226
rect 15967 35266 16007 41186
rect 21927 35266 21967 41186
rect 15967 35226 21967 35266
rect 22338 41186 28338 41226
rect 22338 35266 22378 41186
rect 28298 35266 28338 41186
rect 22338 35226 28338 35266
rect -3146 34815 2854 34855
rect -3146 28895 -3106 34815
rect 2814 28895 2854 34815
rect -3146 28855 2854 28895
rect 3225 34815 9225 34855
rect 3225 28895 3265 34815
rect 9185 28895 9225 34815
rect 3225 28855 9225 28895
rect 9596 34815 15596 34855
rect 9596 28895 9636 34815
rect 15556 28895 15596 34815
rect 9596 28855 15596 28895
rect 15967 34815 21967 34855
rect 15967 28895 16007 34815
rect 21927 28895 21967 34815
rect 15967 28855 21967 28895
rect 22338 34815 28338 34855
rect 22338 28895 22378 34815
rect 28298 28895 28338 34815
rect 22338 28855 28338 28895
rect -3146 28444 2854 28484
rect -3146 22524 -3106 28444
rect 2814 22524 2854 28444
rect -3146 22484 2854 22524
rect 3225 28444 9225 28484
rect 3225 22524 3265 28444
rect 9185 22524 9225 28444
rect 3225 22484 9225 22524
rect 9596 28444 15596 28484
rect 9596 22524 9636 28444
rect 15556 22524 15596 28444
rect 9596 22484 15596 22524
rect 15967 28444 21967 28484
rect 15967 22524 16007 28444
rect 21927 22524 21967 28444
rect 15967 22484 21967 22524
rect 22338 28444 28338 28484
rect 22338 22524 22378 28444
rect 28298 22524 28338 28444
rect 22338 22484 28338 22524
rect -3146 22073 2854 22113
rect -3146 16153 -3106 22073
rect 2814 16153 2854 22073
rect -3146 16113 2854 16153
rect 3225 22073 9225 22113
rect 3225 16153 3265 22073
rect 9185 16153 9225 22073
rect 3225 16113 9225 16153
rect 9596 22073 15596 22113
rect 9596 16153 9636 22073
rect 15556 16153 15596 22073
rect 9596 16113 15596 16153
rect 15967 22073 21967 22113
rect 15967 16153 16007 22073
rect 21927 16153 21967 22073
rect 15967 16113 21967 16153
rect 22338 22073 28338 22113
rect 22338 16153 22378 22073
rect 28298 16153 28338 22073
rect 22338 16113 28338 16153
rect -3146 15702 2854 15742
rect -3146 9782 -3106 15702
rect 2814 9782 2854 15702
rect -3146 9742 2854 9782
rect 3225 15702 9225 15742
rect 3225 9782 3265 15702
rect 9185 9782 9225 15702
rect 3225 9742 9225 9782
rect 9596 15702 15596 15742
rect 9596 9782 9636 15702
rect 15556 9782 15596 15702
rect 9596 9742 15596 9782
rect 15967 15702 21967 15742
rect 15967 9782 16007 15702
rect 21927 9782 21967 15702
rect 15967 9742 21967 9782
rect 22338 15702 28338 15742
rect 22338 9782 22378 15702
rect 28298 9782 28338 15702
rect 22338 9742 28338 9782
rect -3146 9331 2854 9371
rect -3146 3411 -3106 9331
rect 2814 3411 2854 9331
rect -3146 3371 2854 3411
rect 3225 9331 9225 9371
rect 3225 3411 3265 9331
rect 9185 3411 9225 9331
rect 3225 3371 9225 3411
rect 9596 9331 15596 9371
rect 9596 3411 9636 9331
rect 15556 3411 15596 9331
rect 9596 3371 15596 3411
rect 15967 9331 21967 9371
rect 15967 3411 16007 9331
rect 21927 3411 21967 9331
rect 15967 3371 21967 3411
rect 22338 9331 28338 9371
rect 22338 3411 22378 9331
rect 28298 3411 28338 9331
rect 22338 3371 28338 3411
rect -3146 2960 2854 3000
rect -3146 -2960 -3106 2960
rect 2814 -2960 2854 2960
rect -3146 -3000 2854 -2960
rect 3225 2960 9225 3000
rect 3225 -2960 3265 2960
rect 9185 -2960 9225 2960
rect 3225 -3000 9225 -2960
rect 9596 2960 15596 3000
rect 9596 -2960 9636 2960
rect 15556 -2960 15596 2960
rect 9596 -3000 15596 -2960
rect 15967 2960 21967 3000
rect 15967 -2960 16007 2960
rect 21927 -2960 21967 2960
rect 15967 -3000 21967 -2960
rect 22338 2960 28338 3000
rect 22338 -2960 22378 2960
rect 28298 -2960 28338 2960
rect 22338 -3000 28338 -2960
<< mimcapcontact >>
rect -3106 60750 2814 66670
rect 3265 60750 9185 66670
rect 9636 60750 15556 66670
rect 16007 60750 21927 66670
rect 22378 60750 28298 66670
rect -3106 54379 2814 60299
rect 3265 54379 9185 60299
rect 9636 54379 15556 60299
rect 16007 54379 21927 60299
rect 22378 54379 28298 60299
rect -3106 48008 2814 53928
rect 3265 48008 9185 53928
rect 9636 48008 15556 53928
rect 16007 48008 21927 53928
rect 22378 48008 28298 53928
rect -3106 41637 2814 47557
rect 3265 41637 9185 47557
rect 9636 41637 15556 47557
rect 16007 41637 21927 47557
rect 22378 41637 28298 47557
rect -3106 35266 2814 41186
rect 3265 35266 9185 41186
rect 9636 35266 15556 41186
rect 16007 35266 21927 41186
rect 22378 35266 28298 41186
rect -3106 28895 2814 34815
rect 3265 28895 9185 34815
rect 9636 28895 15556 34815
rect 16007 28895 21927 34815
rect 22378 28895 28298 34815
rect -3106 22524 2814 28444
rect 3265 22524 9185 28444
rect 9636 22524 15556 28444
rect 16007 22524 21927 28444
rect 22378 22524 28298 28444
rect -3106 16153 2814 22073
rect 3265 16153 9185 22073
rect 9636 16153 15556 22073
rect 16007 16153 21927 22073
rect 22378 16153 28298 22073
rect -3106 9782 2814 15702
rect 3265 9782 9185 15702
rect 9636 9782 15556 15702
rect 16007 9782 21927 15702
rect 22378 9782 28298 15702
rect -3106 3411 2814 9331
rect 3265 3411 9185 9331
rect 9636 3411 15556 9331
rect 16007 3411 21927 9331
rect 22378 3411 28298 9331
rect -3106 -2960 2814 2960
rect 3265 -2960 9185 2960
rect 9636 -2960 15556 2960
rect 16007 -2960 21927 2960
rect 22378 -2960 28298 2960
<< metal4 >>
rect -3146 66710 -1463 67041
rect 3225 66710 4908 67041
rect 9596 66710 11279 67041
rect 15967 66710 17650 67041
rect 22338 66710 24021 67041
rect -3146 66670 2854 66710
rect -3146 62393 -3106 66670
rect -3186 60750 -3106 62393
rect 2814 62393 2854 66670
rect 3225 66670 9225 66710
rect 3225 62393 3265 66670
rect 2814 60750 3265 62393
rect 9185 62393 9225 66670
rect 9596 66670 15596 66710
rect 9596 62393 9636 66670
rect 9185 60750 9636 62393
rect 15556 62393 15596 66670
rect 15967 66670 21967 66710
rect 15967 62393 16007 66670
rect 15556 60750 16007 62393
rect 21927 62393 21967 66670
rect 22338 66670 28338 66710
rect 22338 62393 22378 66670
rect 21927 60750 22378 62393
rect 28298 62393 28338 66670
rect 28298 60750 28378 62393
rect -3186 60710 28378 60750
rect -3146 60339 -1463 60710
rect 3225 60339 4908 60710
rect 9596 60339 11279 60710
rect 15967 60339 17650 60710
rect 22338 60339 24021 60710
rect -3146 60299 2854 60339
rect -3146 56022 -3106 60299
rect -3186 54379 -3106 56022
rect 2814 56022 2854 60299
rect 3225 60299 9225 60339
rect 3225 56022 3265 60299
rect 2814 54379 3265 56022
rect 9185 56022 9225 60299
rect 9596 60299 15596 60339
rect 9596 56022 9636 60299
rect 9185 54379 9636 56022
rect 15556 56022 15596 60299
rect 15967 60299 21967 60339
rect 15967 56022 16007 60299
rect 15556 54379 16007 56022
rect 21927 56022 21967 60299
rect 22338 60299 28338 60339
rect 22338 56022 22378 60299
rect 21927 54379 22378 56022
rect 28298 56022 28338 60299
rect 28298 54379 28378 56022
rect -3186 54339 28378 54379
rect -3146 53968 -1463 54339
rect 3225 53968 4908 54339
rect 9596 53968 11279 54339
rect 15967 53968 17650 54339
rect 22338 53968 24021 54339
rect -3146 53928 2854 53968
rect -3146 49651 -3106 53928
rect -3186 48008 -3106 49651
rect 2814 49651 2854 53928
rect 3225 53928 9225 53968
rect 3225 49651 3265 53928
rect 2814 48008 3265 49651
rect 9185 49651 9225 53928
rect 9596 53928 15596 53968
rect 9596 49651 9636 53928
rect 9185 48008 9636 49651
rect 15556 49651 15596 53928
rect 15967 53928 21967 53968
rect 15967 49651 16007 53928
rect 15556 48008 16007 49651
rect 21927 49651 21967 53928
rect 22338 53928 28338 53968
rect 22338 49651 22378 53928
rect 21927 48008 22378 49651
rect 28298 49651 28338 53928
rect 28298 48008 28378 49651
rect -3186 47968 28378 48008
rect -3146 47597 -1463 47968
rect 3225 47597 4908 47968
rect 9596 47597 11279 47968
rect 15967 47597 17650 47968
rect 22338 47597 24021 47968
rect -3146 47557 2854 47597
rect -3146 43280 -3106 47557
rect -3186 41637 -3106 43280
rect 2814 43280 2854 47557
rect 3225 47557 9225 47597
rect 3225 43280 3265 47557
rect 2814 41637 3265 43280
rect 9185 43280 9225 47557
rect 9596 47557 15596 47597
rect 9596 43280 9636 47557
rect 9185 41637 9636 43280
rect 15556 43280 15596 47557
rect 15967 47557 21967 47597
rect 15967 43280 16007 47557
rect 15556 41637 16007 43280
rect 21927 43280 21967 47557
rect 22338 47557 28338 47597
rect 22338 43280 22378 47557
rect 21927 41637 22378 43280
rect 28298 43280 28338 47557
rect 28298 41637 28378 43280
rect -3186 41597 28378 41637
rect -3146 41226 -1463 41597
rect 3225 41226 4908 41597
rect 9596 41226 11279 41597
rect 15967 41226 17650 41597
rect 22338 41226 24021 41597
rect -3146 41186 2854 41226
rect -3146 36909 -3106 41186
rect -3186 35266 -3106 36909
rect 2814 36909 2854 41186
rect 3225 41186 9225 41226
rect 3225 36909 3265 41186
rect 2814 35266 3265 36909
rect 9185 36909 9225 41186
rect 9596 41186 15596 41226
rect 9596 36909 9636 41186
rect 9185 35266 9636 36909
rect 15556 36909 15596 41186
rect 15967 41186 21967 41226
rect 15967 36909 16007 41186
rect 15556 35266 16007 36909
rect 21927 36909 21967 41186
rect 22338 41186 28338 41226
rect 22338 36909 22378 41186
rect 21927 35266 22378 36909
rect 28298 36909 28338 41186
rect 28298 35266 28378 36909
rect -3186 35226 28378 35266
rect -3146 34855 -1463 35226
rect 3225 34855 4908 35226
rect 9596 34855 11279 35226
rect 15967 34855 17650 35226
rect 22338 34855 24021 35226
rect -3146 34815 2854 34855
rect -3146 30538 -3106 34815
rect -3186 28895 -3106 30538
rect 2814 30538 2854 34815
rect 3225 34815 9225 34855
rect 3225 30538 3265 34815
rect 2814 28895 3265 30538
rect 9185 30538 9225 34815
rect 9596 34815 15596 34855
rect 9596 30538 9636 34815
rect 9185 28895 9636 30538
rect 15556 30538 15596 34815
rect 15967 34815 21967 34855
rect 15967 30538 16007 34815
rect 15556 28895 16007 30538
rect 21927 30538 21967 34815
rect 22338 34815 28338 34855
rect 22338 30538 22378 34815
rect 21927 28895 22378 30538
rect 28298 30538 28338 34815
rect 28298 28895 28378 30538
rect -3186 28855 28378 28895
rect -3146 28484 -1463 28855
rect 3225 28484 4908 28855
rect 9596 28484 11279 28855
rect 15967 28484 17650 28855
rect 22338 28484 24021 28855
rect -3146 28444 2854 28484
rect -3146 24167 -3106 28444
rect -3186 22524 -3106 24167
rect 2814 24167 2854 28444
rect 3225 28444 9225 28484
rect 3225 24167 3265 28444
rect 2814 22524 3265 24167
rect 9185 24167 9225 28444
rect 9596 28444 15596 28484
rect 9596 24167 9636 28444
rect 9185 22524 9636 24167
rect 15556 24167 15596 28444
rect 15967 28444 21967 28484
rect 15967 24167 16007 28444
rect 15556 22524 16007 24167
rect 21927 24167 21967 28444
rect 22338 28444 28338 28484
rect 22338 24167 22378 28444
rect 21927 22524 22378 24167
rect 28298 24167 28338 28444
rect 28298 22524 28378 24167
rect -3186 22484 28378 22524
rect -3146 22113 -1463 22484
rect 3225 22113 4908 22484
rect 9596 22113 11279 22484
rect 15967 22113 17650 22484
rect 22338 22113 24021 22484
rect -3146 22073 2854 22113
rect -3146 17796 -3106 22073
rect -3186 16153 -3106 17796
rect 2814 17796 2854 22073
rect 3225 22073 9225 22113
rect 3225 17796 3265 22073
rect 2814 16153 3265 17796
rect 9185 17796 9225 22073
rect 9596 22073 15596 22113
rect 9596 17796 9636 22073
rect 9185 16153 9636 17796
rect 15556 17796 15596 22073
rect 15967 22073 21967 22113
rect 15967 17796 16007 22073
rect 15556 16153 16007 17796
rect 21927 17796 21967 22073
rect 22338 22073 28338 22113
rect 22338 17796 22378 22073
rect 21927 16153 22378 17796
rect 28298 17796 28338 22073
rect 28298 16153 28378 17796
rect -3186 16113 28378 16153
rect -3146 15742 -1463 16113
rect 3225 15742 4908 16113
rect 9596 15742 11279 16113
rect 15967 15742 17650 16113
rect 22338 15742 24021 16113
rect -3146 15702 2854 15742
rect -3146 11425 -3106 15702
rect -3186 9782 -3106 11425
rect 2814 11425 2854 15702
rect 3225 15702 9225 15742
rect 3225 11425 3265 15702
rect 2814 9782 3265 11425
rect 9185 11425 9225 15702
rect 9596 15702 15596 15742
rect 9596 11425 9636 15702
rect 9185 9782 9636 11425
rect 15556 11425 15596 15702
rect 15967 15702 21967 15742
rect 15967 11425 16007 15702
rect 15556 9782 16007 11425
rect 21927 11425 21967 15702
rect 22338 15702 28338 15742
rect 22338 11425 22378 15702
rect 21927 9782 22378 11425
rect 28298 11425 28338 15702
rect 28298 9782 28378 11425
rect -3186 9742 28378 9782
rect -3146 9371 -1463 9742
rect 3225 9371 4908 9742
rect 9596 9371 11279 9742
rect 15967 9371 17650 9742
rect 22338 9371 24021 9742
rect -3146 9331 2854 9371
rect -3146 5054 -3106 9331
rect -3186 3411 -3106 5054
rect 2814 5054 2854 9331
rect 3225 9331 9225 9371
rect 3225 5054 3265 9331
rect 2814 3411 3265 5054
rect 9185 5054 9225 9331
rect 9596 9331 15596 9371
rect 9596 5054 9636 9331
rect 9185 3411 9636 5054
rect 15556 5054 15596 9331
rect 15967 9331 21967 9371
rect 15967 5054 16007 9331
rect 15556 3411 16007 5054
rect 21927 5054 21967 9331
rect 22338 9331 28338 9371
rect 22338 5054 22378 9331
rect 21927 3411 22378 5054
rect 28298 5054 28338 9331
rect 28298 3411 28378 5054
rect -3186 3371 28378 3411
rect -3146 3000 -1463 3371
rect 3225 3000 4908 3371
rect 9596 3000 11279 3371
rect 15967 3000 17650 3371
rect 22338 3000 24021 3371
rect -3146 2960 2854 3000
rect -3146 -1317 -3106 2960
rect -3186 -2960 -3106 -1317
rect 2814 -1317 2854 2960
rect 3225 2960 9225 3000
rect 3225 -1317 3265 2960
rect 2814 -2960 3265 -1317
rect 9185 -1317 9225 2960
rect 9596 2960 15596 3000
rect 9596 -1317 9636 2960
rect 9185 -2960 9636 -1317
rect 15556 -1317 15596 2960
rect 15967 2960 21967 3000
rect 15967 -1317 16007 2960
rect 15556 -2960 16007 -1317
rect 21927 -1317 21967 2960
rect 22338 2960 28338 3000
rect 22338 -1317 22378 2960
rect 21927 -2960 22378 -1317
rect 28298 -1317 28338 2960
rect 28298 -2960 28378 -1317
rect -3186 -3000 28378 -2960
rect -3146 -3040 -1463 -3000
rect 3225 -3040 4908 -3000
rect 9596 -3040 11279 -3000
rect 15967 -3040 17650 -3000
rect 22338 -3040 24021 -3000
<< properties >>
string FIXED_BBOX -3186 -3040 2894 3040
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 30 l 30 val 1.822k carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
