magic
tech sky130A
magscale 1 2
timestamp 1658998185
<< nwell >>
rect -358 -288 358 288
<< pmos >>
rect -158 -70 -128 70
rect -62 -70 -32 70
rect 34 -70 64 70
rect 130 -70 160 70
<< pdiff >>
rect -220 58 -158 70
rect -220 -58 -208 58
rect -174 -58 -158 58
rect -220 -70 -158 -58
rect -128 58 -62 70
rect -128 -58 -112 58
rect -78 -58 -62 58
rect -128 -70 -62 -58
rect -32 58 34 70
rect -32 -58 -16 58
rect 18 -58 34 58
rect -32 -70 34 -58
rect 64 58 130 70
rect 64 -58 80 58
rect 114 -58 130 58
rect 64 -70 130 -58
rect 160 58 222 70
rect 160 -58 176 58
rect 210 -58 222 58
rect 160 -70 222 -58
<< pdiffc >>
rect -208 -58 -174 58
rect -112 -58 -78 58
rect -16 -58 18 58
rect 80 -58 114 58
rect 176 -58 210 58
<< nsubdiff >>
rect -322 218 -226 252
rect 226 218 322 252
rect -322 156 -288 218
rect 288 156 322 218
rect -322 -218 -288 -156
rect 288 -218 322 -156
rect -322 -252 -226 -218
rect 226 -252 322 -218
<< nsubdiffcont >>
rect -226 218 226 252
rect -322 -156 -288 156
rect 288 -156 322 156
rect -226 -252 226 -218
<< poly >>
rect -80 151 82 167
rect -80 117 -64 151
rect -30 117 32 151
rect 66 117 82 151
rect -80 101 82 117
rect -158 70 -128 96
rect -62 70 -32 101
rect 34 70 64 101
rect 130 70 160 96
rect -158 -101 -128 -70
rect -62 -96 -32 -70
rect 34 -96 64 -70
rect 130 -101 160 -70
rect -176 -117 -110 -101
rect -176 -151 -160 -117
rect -126 -151 -110 -117
rect -176 -167 -110 -151
rect 112 -117 178 -101
rect 112 -151 128 -117
rect 162 -151 178 -117
rect 112 -167 178 -151
<< polycont >>
rect -64 117 -30 151
rect 32 117 66 151
rect -160 -151 -126 -117
rect 128 -151 162 -117
<< locali >>
rect -322 218 -226 252
rect 226 218 322 252
rect -322 156 -288 218
rect 288 156 322 218
rect -80 117 -64 151
rect -30 117 32 151
rect 66 117 82 151
rect -208 58 -174 74
rect -208 -74 -174 -58
rect -112 58 -78 74
rect -112 -74 -78 -58
rect -16 58 18 74
rect -16 -74 18 -58
rect 80 58 114 74
rect 80 -74 114 -58
rect 176 58 210 74
rect 176 -74 210 -58
rect -176 -151 -160 -117
rect -126 -151 -110 -117
rect 112 -151 128 -117
rect 162 -151 178 -117
rect -322 -218 -288 -156
rect 288 -218 322 -156
rect -322 -252 -226 -218
rect 226 -252 322 -218
<< viali >>
rect -64 117 -30 151
rect 32 117 66 151
rect -208 -58 -174 58
rect -112 -58 -78 58
rect -16 -58 18 58
rect 80 -58 114 58
rect 176 -58 210 58
rect -160 -151 -126 -117
rect 128 -151 162 -117
<< metal1 >>
rect -64 157 -30 288
rect -76 151 -18 157
rect 20 151 78 157
rect -76 117 -64 151
rect -30 117 32 151
rect 66 117 78 151
rect -76 111 -18 117
rect 20 111 78 117
rect -224 58 -158 70
rect -224 -58 -218 58
rect -166 -58 -158 58
rect -224 -70 -158 -58
rect -128 58 -62 70
rect -128 -58 -122 58
rect -70 -58 -62 58
rect -128 -70 -62 -58
rect -32 58 34 70
rect -32 -58 -26 58
rect 26 -58 34 58
rect -32 -70 34 -58
rect 64 58 130 70
rect 64 -58 70 58
rect 124 -58 130 58
rect 64 -70 130 -58
rect 160 58 226 70
rect 160 -58 166 58
rect 220 -58 226 58
rect 160 -70 226 -58
rect -172 -117 -114 -111
rect 116 -117 174 -111
rect -172 -151 -160 -117
rect -126 -151 128 -117
rect 162 -151 174 -117
rect -172 -157 -114 -151
rect 116 -157 174 -151
<< via1 >>
rect -218 -58 -208 58
rect -208 -58 -174 58
rect -174 -58 -166 58
rect -122 -58 -112 58
rect -112 -58 -78 58
rect -78 -58 -70 58
rect -26 -58 -16 58
rect -16 -58 18 58
rect 18 -58 26 58
rect 70 -58 80 58
rect 80 -58 114 58
rect 114 -58 124 58
rect 166 -58 176 58
rect 176 -58 210 58
rect 210 -58 220 58
<< metal2 >>
rect -16 70 18 288
rect -225 58 -158 70
rect -225 -58 -220 58
rect -164 -58 -158 58
rect -225 -70 -158 -58
rect -128 58 -62 70
rect -128 -58 -124 58
rect -68 -58 -62 58
rect -128 -70 -62 -58
rect -32 58 34 70
rect -32 -58 -26 58
rect 26 -58 34 58
rect -32 -70 34 -58
rect 64 58 130 70
rect 64 -58 70 58
rect 126 -58 130 58
rect 64 -70 130 -58
rect 160 58 227 70
rect 160 -58 166 58
rect 222 -58 227 58
rect 160 -70 227 -58
<< via2 >>
rect -220 -58 -218 58
rect -218 -58 -166 58
rect -166 -58 -164 58
rect -124 -58 -122 58
rect -122 -58 -70 58
rect -70 -58 -68 58
rect 70 -58 124 58
rect 124 -58 126 58
rect 166 -58 220 58
rect 220 -58 222 58
<< metal3 >>
rect -225 58 -62 70
rect -225 -58 -220 58
rect -164 -58 -124 58
rect -68 -10 -62 58
rect 64 58 227 70
rect 64 -10 70 58
rect -68 -58 70 -10
rect 126 -58 166 58
rect 222 -58 227 58
rect -225 -70 227 -58
<< properties >>
string FIXED_BBOX -306 -236 306 236
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.7 l 0.15 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
