magic
tech sky130A
magscale 1 2
timestamp 1668357910
<< pwell >>
rect -455 -280 455 280
<< nmoslvt >>
rect -255 -70 -225 70
rect -159 -70 -129 70
rect -63 -70 -33 70
rect 33 -70 63 70
rect 129 -70 159 70
rect 225 -70 255 70
<< ndiff >>
rect -317 58 -255 70
rect -317 -58 -305 58
rect -271 -58 -255 58
rect -317 -70 -255 -58
rect -225 58 -159 70
rect -225 -58 -209 58
rect -175 -58 -159 58
rect -225 -70 -159 -58
rect -129 58 -63 70
rect -129 -58 -113 58
rect -79 -58 -63 58
rect -129 -70 -63 -58
rect -33 58 33 70
rect -33 -58 -17 58
rect 17 -58 33 58
rect -33 -70 33 -58
rect 63 58 129 70
rect 63 -58 79 58
rect 113 -58 129 58
rect 63 -70 129 -58
rect 159 58 225 70
rect 159 -58 175 58
rect 209 -58 225 58
rect 159 -70 225 -58
rect 255 58 317 70
rect 255 -58 271 58
rect 305 -58 317 58
rect 255 -70 317 -58
<< ndiffc >>
rect -305 -58 -271 58
rect -209 -58 -175 58
rect -113 -58 -79 58
rect -17 -58 17 58
rect 79 -58 113 58
rect 175 -58 209 58
rect 271 -58 305 58
<< psubdiff >>
rect -419 210 -323 244
rect 323 210 419 244
rect -419 148 -385 210
rect 385 148 419 210
rect -419 -210 -385 -148
rect 385 -210 419 -148
rect -419 -244 -323 -210
rect 323 -244 419 -210
<< psubdiffcont >>
rect -323 210 323 244
rect -419 -148 -385 148
rect 385 -148 419 148
rect -323 -244 323 -210
<< poly >>
rect -273 142 -207 158
rect -273 108 -257 142
rect -223 108 -207 142
rect -273 92 -207 108
rect 207 142 273 158
rect 207 108 223 142
rect 257 108 273 142
rect -255 70 -225 92
rect -159 70 -129 96
rect -63 70 -33 96
rect 33 70 63 97
rect 129 70 159 96
rect 207 92 273 108
rect 225 70 255 92
rect -255 -97 -225 -70
rect -159 -92 -129 -70
rect -63 -92 -33 -70
rect -177 -108 -33 -92
rect -177 -142 -161 -108
rect -127 -142 -33 -108
rect -177 -158 -33 -142
rect 33 -92 63 -70
rect 129 -92 159 -70
rect 33 -108 177 -92
rect 225 -96 255 -70
rect 33 -142 127 -108
rect 161 -142 177 -108
rect 33 -158 177 -142
<< polycont >>
rect -257 108 -223 142
rect 223 108 257 142
rect -161 -142 -127 -108
rect 127 -142 161 -108
<< locali >>
rect -419 210 -323 244
rect 323 210 419 244
rect -419 148 -385 210
rect 385 148 419 210
rect -273 108 -257 142
rect -223 108 -207 142
rect 207 108 223 142
rect 257 108 273 142
rect -305 58 -271 74
rect -305 -74 -271 -58
rect -209 58 -175 74
rect -209 -74 -175 -58
rect -113 58 -79 74
rect -113 -74 -79 -58
rect -17 58 17 74
rect -17 -74 17 -58
rect 79 58 113 74
rect 79 -74 113 -58
rect 175 58 209 74
rect 175 -74 209 -58
rect 271 58 305 74
rect 271 -74 305 -58
rect -177 -142 -161 -108
rect -127 -142 -111 -108
rect 111 -142 127 -108
rect 161 -142 177 -108
rect -419 -210 -385 -148
rect 385 -210 419 -148
rect -419 -244 -323 -210
rect 323 -244 419 -210
<< viali >>
rect -257 108 -223 142
rect 223 108 257 142
rect -305 -58 -271 58
rect -209 -58 -175 58
rect -113 -58 -79 57
rect -17 -58 17 58
rect 79 -58 113 58
rect 175 -58 209 58
rect 271 -58 305 58
rect -161 -142 -127 -108
rect 127 -142 161 -108
<< metal1 >>
rect -305 142 -211 148
rect -305 108 -257 142
rect -223 108 -211 142
rect -305 102 -211 108
rect -305 70 -269 102
rect -113 70 -79 279
rect 79 70 113 280
rect 211 142 305 148
rect 211 108 223 142
rect 257 108 305 142
rect 211 102 305 108
rect 269 70 305 102
rect -318 58 -162 70
rect -318 -58 -314 58
rect -262 -58 -218 58
rect -166 -58 -162 58
rect -318 -70 -162 -58
rect -119 57 -73 70
rect -119 -58 -113 57
rect -79 -58 -73 57
rect -119 -70 -73 -58
rect -30 58 30 70
rect -30 -58 -26 58
rect 26 -58 30 58
rect -30 -70 30 -58
rect 73 58 119 70
rect 73 -58 79 58
rect 113 -58 119 58
rect 73 -70 119 -58
rect 162 58 318 70
rect 162 -58 166 58
rect 218 -58 262 58
rect 314 -58 318 58
rect 162 -70 318 -58
rect -173 -108 -115 -102
rect -455 -142 -161 -108
rect -127 -142 -115 -108
rect -173 -148 -115 -142
rect 115 -108 173 -102
rect 115 -142 127 -108
rect 161 -142 455 -108
rect 115 -148 173 -142
<< via1 >>
rect -314 -58 -305 58
rect -305 -58 -271 58
rect -271 -58 -262 58
rect -218 -58 -209 58
rect -209 -58 -175 58
rect -175 -58 -166 58
rect -26 -58 -17 58
rect -17 -58 17 58
rect 17 -58 26 58
rect 166 -58 175 58
rect 175 -58 209 58
rect 209 -58 218 58
rect 262 -58 271 58
rect 271 -58 305 58
rect 305 -58 314 58
<< metal2 >>
rect -318 58 -162 70
rect -318 -58 -314 58
rect -262 -58 -218 58
rect -166 -10 -162 58
rect -30 58 30 70
rect -30 -10 -26 58
rect -166 -58 -26 -10
rect 26 -10 30 58
rect 162 58 318 70
rect 162 -10 166 58
rect 26 -58 166 -10
rect 218 -58 262 58
rect 314 -58 318 58
rect -318 -70 318 -58
<< properties >>
string FIXED_BBOX -402 -227 402 227
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 0.7 l 0.150 m 1 nf 6 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
