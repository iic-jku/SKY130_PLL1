magic
tech sky130A
magscale 1 2
timestamp 1666523630
<< nwell >>
rect -647 -289 647 289
<< pmos >>
rect -447 -70 -417 70
rect -351 -70 -321 70
rect -255 -70 -225 70
rect -159 -70 -129 70
rect -63 -70 -33 70
rect 33 -70 63 70
rect 129 -70 159 70
rect 225 -70 255 70
rect 321 -70 351 70
rect 417 -70 447 70
<< pdiff >>
rect -509 58 -447 70
rect -509 -58 -497 58
rect -463 -58 -447 58
rect -509 -70 -447 -58
rect -417 58 -351 70
rect -417 -58 -401 58
rect -367 -58 -351 58
rect -417 -70 -351 -58
rect -321 58 -255 70
rect -321 -58 -305 58
rect -271 -58 -255 58
rect -321 -70 -255 -58
rect -225 58 -159 70
rect -225 -58 -209 58
rect -175 -58 -159 58
rect -225 -70 -159 -58
rect -129 58 -63 70
rect -129 -58 -113 58
rect -79 -58 -63 58
rect -129 -70 -63 -58
rect -33 58 33 70
rect -33 -58 -17 58
rect 17 -58 33 58
rect -33 -70 33 -58
rect 63 58 129 70
rect 63 -58 79 58
rect 113 -58 129 58
rect 63 -70 129 -58
rect 159 58 225 70
rect 159 -58 175 58
rect 209 -58 225 58
rect 159 -70 225 -58
rect 255 58 321 70
rect 255 -58 271 58
rect 305 -58 321 58
rect 255 -70 321 -58
rect 351 58 417 70
rect 351 -58 367 58
rect 401 -58 417 58
rect 351 -70 417 -58
rect 447 58 510 70
rect 447 -58 463 58
rect 497 0 510 58
rect 497 -58 509 0
rect 447 -70 509 -58
<< pdiffc >>
rect -497 -58 -463 58
rect -401 -58 -367 58
rect -305 -58 -271 58
rect -209 -58 -175 58
rect -113 -58 -79 58
rect -17 -58 17 58
rect 79 -58 113 58
rect 175 -58 209 58
rect 271 -58 305 58
rect 367 -58 401 58
rect 463 -58 497 58
<< nsubdiff >>
rect -611 219 -515 253
rect 515 219 611 253
rect -611 157 -577 219
rect 577 157 611 219
rect -611 -219 -577 -157
rect 577 -219 611 -157
rect -611 -253 -515 -219
rect 515 -253 611 -219
<< nsubdiffcont >>
rect -515 219 515 253
rect -611 -157 -577 157
rect 577 -157 611 157
rect -515 -253 515 -219
<< poly >>
rect -465 151 -399 167
rect -465 117 -449 151
rect -415 117 -399 151
rect -465 101 -399 117
rect 399 151 465 167
rect 399 117 415 151
rect 449 117 465 151
rect 399 101 465 117
rect -447 70 -417 101
rect -351 70 -321 96
rect -255 70 -225 96
rect -159 70 -129 96
rect -63 70 -33 96
rect 33 70 63 96
rect 129 70 159 96
rect 225 70 255 96
rect 321 70 351 96
rect 417 70 447 101
rect -447 -96 -417 -70
rect -351 -101 -321 -70
rect -255 -101 -225 -70
rect -159 -101 -129 -70
rect -63 -101 -33 -70
rect 33 -101 63 -70
rect 129 -101 159 -70
rect 225 -101 255 -70
rect 321 -101 351 -70
rect 417 -96 447 -70
rect -369 -117 369 -101
rect -369 -151 -353 -117
rect -319 -151 -257 -117
rect -223 -151 -161 -117
rect -127 -151 -65 -117
rect -31 -151 31 -117
rect 65 -151 127 -117
rect 161 -151 223 -117
rect 257 -151 319 -117
rect 353 -151 369 -117
rect -369 -167 369 -151
<< polycont >>
rect -449 117 -415 151
rect 415 117 449 151
rect -353 -151 -319 -117
rect -257 -151 -223 -117
rect -161 -151 -127 -117
rect -65 -151 -31 -117
rect 31 -151 65 -117
rect 127 -151 161 -117
rect 223 -151 257 -117
rect 319 -151 353 -117
<< locali >>
rect -611 219 -515 253
rect 515 219 611 253
rect -611 157 -577 219
rect 577 157 611 219
rect -465 117 -449 151
rect -415 117 -399 151
rect 399 117 415 151
rect 449 117 465 151
rect -497 58 -463 74
rect -497 -74 -463 -58
rect -401 58 -367 74
rect -401 -74 -367 -58
rect -305 58 -271 74
rect -305 -74 -271 -58
rect -209 58 -175 74
rect -209 -74 -175 -58
rect -113 58 -79 74
rect -113 -74 -79 -58
rect -17 58 17 74
rect -17 -74 17 -58
rect 79 58 113 74
rect 79 -74 113 -58
rect 175 58 209 74
rect 175 -74 209 -58
rect 271 58 305 74
rect 271 -74 305 -58
rect 367 58 401 74
rect 367 -74 401 -58
rect 463 58 497 74
rect 463 -74 497 -58
rect -369 -151 -353 -117
rect -319 -151 -257 -117
rect -223 -151 -161 -117
rect -127 -151 -65 -117
rect -31 -151 31 -117
rect 65 -151 127 -117
rect 161 -151 223 -117
rect 257 -151 319 -117
rect 353 -151 369 -117
rect -611 -219 -577 -157
rect 577 -219 611 -157
rect -611 -253 -515 -219
rect 515 -253 611 -219
<< viali >>
rect -449 117 -415 151
rect 415 117 449 151
rect -497 -58 -463 58
rect -401 -58 -367 58
rect -305 -58 -271 58
rect -209 -58 -175 58
rect -113 -58 -79 58
rect -17 -58 17 58
rect 79 -58 113 58
rect 175 -58 209 58
rect 271 -58 305 58
rect 367 -58 401 58
rect 463 -58 497 58
rect -353 -151 -319 -117
rect -257 -151 -223 -117
rect -161 -151 -127 -117
rect -65 -151 -31 -117
rect 31 -151 65 -117
rect 127 -151 161 -117
rect 223 -151 257 -117
rect 319 -151 353 -117
<< metal1 >>
rect -461 151 -403 157
rect 403 151 461 157
rect -461 117 -449 151
rect -415 117 415 151
rect 449 117 461 151
rect -461 111 -403 117
rect 403 111 461 117
rect -508 60 -354 70
rect -508 8 -505 60
rect -453 8 -409 60
rect -357 8 -354 60
rect -508 0 -497 8
rect -503 -58 -497 0
rect -463 0 -401 8
rect -463 -58 -457 0
rect -503 -70 -457 -58
rect -407 -58 -401 0
rect -367 0 -354 8
rect -311 58 -265 70
rect -311 0 -305 58
rect -367 -58 -361 0
rect -407 -70 -361 -58
rect -317 -8 -305 0
rect -271 0 -265 58
rect -220 60 -162 70
rect -220 8 -217 60
rect -165 8 -162 60
rect -220 0 -209 8
rect -271 -8 -259 0
rect -317 -60 -314 -8
rect -262 -60 -259 -8
rect -317 -70 -259 -60
rect -215 -58 -209 0
rect -175 0 -162 8
rect -119 58 -73 70
rect -119 0 -113 58
rect -175 -58 -169 0
rect -215 -70 -169 -58
rect -125 -8 -113 0
rect -79 0 -73 58
rect -28 60 30 70
rect -28 8 -25 60
rect 27 8 30 60
rect -28 0 -17 8
rect -79 -8 -67 0
rect -125 -60 -122 -8
rect -70 -60 -67 -8
rect -125 -70 -67 -60
rect -23 -58 -17 0
rect 17 0 30 8
rect 73 58 119 70
rect 73 0 79 58
rect 17 -58 23 0
rect -23 -70 23 -58
rect 67 -8 79 0
rect 113 0 119 58
rect 164 60 222 70
rect 164 8 167 60
rect 219 8 222 60
rect 164 0 175 8
rect 113 -8 125 0
rect 67 -60 70 -8
rect 122 -60 125 -8
rect 67 -70 125 -60
rect 169 -58 175 0
rect 209 0 222 8
rect 265 58 311 70
rect 265 0 271 58
rect 209 -58 215 0
rect 169 -70 215 -58
rect 259 -8 271 0
rect 305 0 311 58
rect 356 60 510 70
rect 356 8 359 60
rect 411 8 455 60
rect 507 8 510 60
rect 356 0 367 8
rect 305 -8 317 0
rect 259 -60 262 -8
rect 314 -60 317 -8
rect 259 -70 317 -60
rect 361 -58 367 0
rect 401 0 463 8
rect 401 -58 407 0
rect 361 -70 407 -58
rect 457 -58 463 0
rect 497 0 510 8
rect 497 -58 503 0
rect 457 -70 503 -58
rect -365 -117 365 -111
rect -365 -151 -353 -117
rect -319 -151 -257 -117
rect -223 -151 -161 -117
rect -127 -151 -65 -117
rect -31 -151 31 -117
rect 65 -151 127 -117
rect 161 -151 223 -117
rect 257 -151 319 -117
rect 353 -151 365 -117
rect -365 -157 365 -151
<< via1 >>
rect -505 58 -453 60
rect -505 8 -497 58
rect -497 8 -463 58
rect -463 8 -453 58
rect -409 58 -357 60
rect -409 8 -401 58
rect -401 8 -367 58
rect -367 8 -357 58
rect -217 58 -165 60
rect -217 8 -209 58
rect -209 8 -175 58
rect -175 8 -165 58
rect -314 -58 -305 -8
rect -305 -58 -271 -8
rect -271 -58 -262 -8
rect -314 -60 -262 -58
rect -25 58 27 60
rect -25 8 -17 58
rect -17 8 17 58
rect 17 8 27 58
rect -122 -58 -113 -8
rect -113 -58 -79 -8
rect -79 -58 -70 -8
rect -122 -60 -70 -58
rect 167 58 219 60
rect 167 8 175 58
rect 175 8 209 58
rect 209 8 219 58
rect 70 -58 79 -8
rect 79 -58 113 -8
rect 113 -58 122 -8
rect 70 -60 122 -58
rect 359 58 411 60
rect 359 8 367 58
rect 367 8 401 58
rect 401 8 411 58
rect 455 58 507 60
rect 455 8 463 58
rect 463 8 497 58
rect 497 8 507 58
rect 262 -58 271 -8
rect 271 -58 305 -8
rect 305 -58 314 -8
rect 262 -60 314 -58
<< metal2 >>
rect -508 60 510 70
rect -508 8 -505 60
rect -453 8 -409 60
rect -357 28 -217 60
rect -357 8 -354 28
rect -508 0 -354 8
rect -220 8 -217 28
rect -165 28 -25 60
rect -165 8 -162 28
rect -220 0 -162 8
rect -28 8 -25 28
rect 27 28 167 60
rect 27 8 30 28
rect -28 0 30 8
rect 164 8 167 28
rect 219 28 359 60
rect 219 8 222 28
rect 164 0 222 8
rect 356 8 359 28
rect 411 8 455 60
rect 507 8 510 60
rect 356 0 510 8
rect -317 -8 -259 0
rect -317 -60 -314 -8
rect -262 -28 -259 -8
rect -125 -8 -67 0
rect -125 -28 -122 -8
rect -262 -60 -122 -28
rect -70 -28 -67 -8
rect 67 -8 125 0
rect 67 -28 70 -8
rect -70 -60 70 -28
rect 122 -28 125 -8
rect 259 -8 317 0
rect 259 -28 262 -8
rect 122 -60 262 -28
rect 314 -60 317 -8
rect -317 -70 317 -60
<< properties >>
string FIXED_BBOX -594 -236 594 236
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.7 l 0.15 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
