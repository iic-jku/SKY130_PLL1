magic
tech sky130A
timestamp 1668153059
<< metal3 >>
rect -325 -300 275 300
<< mimcap >>
rect -275 230 225 250
rect -275 -230 -255 230
rect 205 -230 225 230
rect -275 -250 225 -230
<< mimcapcontact >>
rect -255 -230 205 230
<< metal4 >>
rect -275 230 225 250
rect -275 -230 -255 230
rect 205 -230 225 230
rect -275 -250 225 -230
<< properties >>
string FIXED_BBOX -325 -300 275 300
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 5 l 5 val 53.8 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
