magic
tech sky130A
magscale 1 2
timestamp 1654967793
<< error_p >>
rect -365 -108 -307 -102
rect 307 -108 365 -102
rect -365 -142 -353 -108
rect 307 -142 319 -108
rect -365 -148 -307 -142
rect 307 -148 365 -142
<< pwell >>
rect -551 -280 551 280
<< nmos >>
rect -351 -70 -321 70
rect -255 -70 -225 70
rect -159 -70 -129 70
rect -63 -70 -33 70
rect 33 -70 63 70
rect 129 -70 159 70
rect 225 -70 255 70
rect 321 -70 351 70
<< ndiff >>
rect -413 58 -351 70
rect -413 -58 -401 58
rect -367 -58 -351 58
rect -413 -70 -351 -58
rect -321 58 -255 70
rect -321 -58 -305 58
rect -271 -58 -255 58
rect -321 -70 -255 -58
rect -225 58 -159 70
rect -225 -58 -209 58
rect -175 -58 -159 58
rect -225 -70 -159 -58
rect -129 58 -63 70
rect -129 -58 -113 58
rect -79 -58 -63 58
rect -129 -70 -63 -58
rect -33 58 33 70
rect -33 -58 -17 58
rect 17 -58 33 58
rect -33 -70 33 -58
rect 63 58 129 70
rect 63 -58 79 58
rect 113 -58 129 58
rect 63 -70 129 -58
rect 159 58 225 70
rect 159 -58 175 58
rect 209 -58 225 58
rect 159 -70 225 -58
rect 255 58 321 70
rect 255 -58 271 58
rect 305 -58 321 58
rect 255 -70 321 -58
rect 351 58 413 70
rect 351 -58 367 58
rect 401 -58 413 58
rect 351 -70 413 -58
<< ndiffc >>
rect -401 -58 -367 58
rect -305 -58 -271 58
rect -209 -58 -175 58
rect -113 -58 -79 58
rect -17 -58 17 58
rect 79 -58 113 58
rect 175 -58 209 58
rect 271 -58 305 58
rect 367 -58 401 58
<< psubdiff >>
rect -515 210 -419 244
rect 419 210 515 244
rect -515 148 -481 210
rect 481 148 515 210
rect -515 -210 -481 -148
rect 481 -210 515 -148
rect -515 -244 -419 -210
rect 419 -244 515 -210
<< psubdiffcont >>
rect -419 210 419 244
rect -515 -148 -481 148
rect 481 -148 515 148
rect -419 -244 419 -210
<< poly >>
rect -273 142 -111 158
rect -273 108 -257 142
rect -223 108 -161 142
rect -127 108 -111 142
rect -351 70 -321 96
rect -273 92 -111 108
rect 111 142 273 158
rect 111 108 127 142
rect 161 108 223 142
rect 257 108 273 142
rect -255 70 -225 92
rect -159 70 -129 92
rect -63 70 -33 96
rect 33 70 63 96
rect 111 92 273 108
rect 129 70 159 92
rect 225 70 255 92
rect 321 70 351 96
rect -351 -92 -321 -70
rect -369 -108 -303 -92
rect -255 -96 -225 -70
rect -159 -96 -129 -70
rect -63 -92 -33 -70
rect 33 -92 63 -70
rect -369 -142 -353 -108
rect -319 -142 -303 -108
rect -369 -158 -303 -142
rect -81 -108 81 -92
rect 129 -96 159 -70
rect 225 -96 255 -70
rect 321 -92 351 -70
rect -81 -142 -65 -108
rect -31 -142 31 -108
rect 65 -142 81 -108
rect -81 -158 81 -142
rect 303 -108 369 -92
rect 303 -142 319 -108
rect 353 -142 369 -108
rect 303 -158 369 -142
<< polycont >>
rect -257 108 -223 142
rect -161 108 -127 142
rect 127 108 161 142
rect 223 108 257 142
rect -353 -142 -319 -108
rect -65 -142 -31 -108
rect 31 -142 65 -108
rect 319 -142 353 -108
<< locali >>
rect -515 210 -419 244
rect 419 210 515 244
rect -515 148 -481 210
rect 481 148 515 210
rect -273 108 -257 142
rect -223 108 -161 142
rect -127 108 -111 142
rect 111 108 127 142
rect 161 108 223 142
rect 257 108 273 142
rect -401 58 -367 74
rect -401 -74 -367 -58
rect -305 58 -271 74
rect -305 -74 -271 -58
rect -209 58 -175 74
rect -209 -74 -175 -58
rect -113 58 -79 74
rect -113 -74 -79 -58
rect -17 58 17 74
rect -17 -74 17 -58
rect 79 58 113 74
rect 79 -74 113 -58
rect 175 58 209 74
rect 175 -74 209 -58
rect 271 58 305 74
rect 271 -74 305 -58
rect 367 58 401 74
rect 367 -74 401 -58
rect -369 -142 -353 -108
rect -319 -142 -303 -108
rect -81 -142 -65 -108
rect -31 -142 31 -108
rect 65 -142 81 -108
rect 303 -142 319 -108
rect 353 -142 369 -108
rect -515 -210 -481 -148
rect 481 -210 515 -148
rect -515 -244 -419 -210
rect 419 -244 515 -210
<< viali >>
rect -257 108 -223 142
rect -161 108 -127 142
rect 127 108 161 142
rect 223 108 257 142
rect -401 -58 -367 58
rect -305 -58 -271 58
rect -209 -58 -175 58
rect -113 -58 -79 58
rect -17 -58 17 58
rect 79 -58 113 58
rect 175 -58 209 58
rect 271 -58 305 58
rect 367 -58 401 58
rect -353 -142 -319 -108
rect -65 -142 -31 -108
rect 31 -142 65 -108
rect 319 -142 353 -108
<< metal1 >>
rect -269 142 -211 148
rect -173 142 -115 148
rect -269 108 -257 142
rect -223 108 -161 142
rect -127 108 -115 142
rect -269 102 -211 108
rect -173 102 -115 108
rect 115 142 173 148
rect 211 142 269 148
rect 115 108 127 142
rect 161 108 223 142
rect 257 108 269 142
rect 115 102 173 108
rect 211 102 269 108
rect -416 66 -352 70
rect -416 14 -410 66
rect -358 14 -352 66
rect -416 6 -401 14
rect -407 -58 -401 6
rect -367 6 -352 14
rect -320 66 -256 70
rect -320 14 -314 66
rect -262 14 -256 66
rect -320 6 -305 14
rect -367 -58 -361 6
rect -407 -70 -361 -58
rect -311 -58 -305 6
rect -271 6 -256 14
rect -215 58 -169 70
rect -271 -58 -265 6
rect -215 -6 -209 58
rect -311 -70 -265 -58
rect -224 -12 -209 -6
rect -175 -6 -169 58
rect -128 66 -64 70
rect -128 14 -122 66
rect -70 14 -64 66
rect -128 6 -113 14
rect -175 -12 -160 -6
rect -224 -64 -218 -12
rect -166 -64 -160 -12
rect -224 -70 -160 -64
rect -119 -58 -113 6
rect -79 6 -64 14
rect -23 58 23 70
rect -79 -58 -73 6
rect -23 -6 -17 58
rect -119 -70 -73 -58
rect -32 -12 -17 -6
rect 17 -6 23 58
rect 64 66 128 70
rect 64 14 70 66
rect 122 14 128 66
rect 64 6 79 14
rect 17 -12 32 -6
rect -32 -64 -26 -12
rect 26 -64 32 -12
rect -32 -70 32 -64
rect 73 -58 79 6
rect 113 6 128 14
rect 169 58 215 70
rect 113 -58 119 6
rect 169 -6 175 58
rect 73 -70 119 -58
rect 160 -12 175 -6
rect 209 -6 215 58
rect 256 66 320 70
rect 256 14 262 66
rect 314 14 320 66
rect 256 6 271 14
rect 209 -12 224 -6
rect 160 -64 166 -12
rect 218 -64 224 -12
rect 160 -70 224 -64
rect 265 -58 271 6
rect 305 6 320 14
rect 352 66 416 70
rect 352 14 358 66
rect 410 14 416 66
rect 352 6 367 14
rect 305 -58 311 6
rect 265 -70 311 -58
rect 361 -58 367 6
rect 401 6 416 14
rect 401 -58 407 6
rect 361 -70 407 -58
rect -365 -108 -307 -102
rect -365 -142 -353 -108
rect -319 -142 -307 -108
rect -365 -148 -307 -142
rect -77 -108 -19 -102
rect 19 -108 77 -102
rect -77 -142 -65 -108
rect -31 -142 31 -108
rect 65 -142 77 -108
rect -77 -148 -19 -142
rect 19 -148 77 -142
rect 307 -108 365 -102
rect 307 -142 319 -108
rect 353 -142 365 -108
rect 307 -148 365 -142
<< via1 >>
rect -410 58 -358 66
rect -410 14 -401 58
rect -401 14 -367 58
rect -367 14 -358 58
rect -314 58 -262 66
rect -314 14 -305 58
rect -305 14 -271 58
rect -271 14 -262 58
rect -122 58 -70 66
rect -122 14 -113 58
rect -113 14 -79 58
rect -79 14 -70 58
rect -218 -58 -209 -12
rect -209 -58 -175 -12
rect -175 -58 -166 -12
rect -218 -64 -166 -58
rect 70 58 122 66
rect 70 14 79 58
rect 79 14 113 58
rect 113 14 122 58
rect -26 -58 -17 -12
rect -17 -58 17 -12
rect 17 -58 26 -12
rect -26 -64 26 -58
rect 262 58 314 66
rect 262 14 271 58
rect 271 14 305 58
rect 305 14 314 58
rect 166 -58 175 -12
rect 175 -58 209 -12
rect 209 -58 218 -12
rect 166 -64 218 -58
rect 358 58 410 66
rect 358 14 367 58
rect 367 14 401 58
rect 401 14 410 58
<< metal2 >>
rect -421 68 -251 77
rect -421 12 -412 68
rect -356 12 -316 68
rect -260 12 -251 68
rect -421 3 -251 12
rect -133 68 -59 77
rect -133 12 -124 68
rect -68 12 -59 68
rect -133 3 -59 12
rect 59 68 133 77
rect 59 12 68 68
rect 124 12 133 68
rect 59 3 133 12
rect 251 68 421 77
rect 251 12 260 68
rect 316 12 356 68
rect 412 12 421 68
rect 251 3 421 12
rect -224 -12 -160 -6
rect -224 -64 -218 -12
rect -166 -64 -160 -12
rect -224 -70 -160 -64
rect -32 -12 32 -6
rect -32 -64 -26 -12
rect 26 -64 32 -12
rect -32 -70 32 -64
rect 160 -12 224 -6
rect 160 -64 166 -12
rect 218 -64 224 -12
rect 160 -70 224 -64
<< via2 >>
rect -412 66 -356 68
rect -412 14 -410 66
rect -410 14 -358 66
rect -358 14 -356 66
rect -412 12 -356 14
rect -316 66 -260 68
rect -316 14 -314 66
rect -314 14 -262 66
rect -262 14 -260 66
rect -316 12 -260 14
rect -124 66 -68 68
rect -124 14 -122 66
rect -122 14 -70 66
rect -70 14 -68 66
rect -124 12 -68 14
rect 68 66 124 68
rect 68 14 70 66
rect 70 14 122 66
rect 122 14 124 66
rect 68 12 124 14
rect 260 66 316 68
rect 260 14 262 66
rect 262 14 314 66
rect 314 14 316 66
rect 260 12 316 14
rect 356 66 412 68
rect 356 14 358 66
rect 358 14 410 66
rect 410 14 412 66
rect 356 12 412 14
<< metal3 >>
rect -421 70 -251 77
rect -133 70 -59 77
rect 59 70 133 77
rect 251 70 421 77
rect -421 68 421 70
rect -421 12 -412 68
rect -356 12 -316 68
rect -260 12 -124 68
rect -68 12 68 68
rect 124 12 260 68
rect 316 12 356 68
rect 412 12 421 68
rect -421 10 421 12
rect -421 3 -251 10
rect -133 3 -59 10
rect 59 3 133 10
rect 251 3 421 10
<< properties >>
string FIXED_BBOX -498 -227 498 227
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.7 l 0.150 m 1 nf 8 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
