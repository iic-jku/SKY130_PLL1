magic
tech sky130A
magscale 1 2
timestamp 1668357910
<< metal2 >>
rect 73442 12503 74458 12600
rect 73440 12331 74458 12503
rect 71224 10791 71794 11361
rect 73440 11215 73658 12331
rect 74253 11215 74458 12331
rect 73440 10942 74458 11215
rect 69774 6219 70206 6651
<< via2 >>
rect 73658 11215 74253 12331
<< metal3 >>
rect 73440 12331 74458 19661
rect 73440 11215 73658 12331
rect 74253 11215 74458 12331
rect 73440 10942 74458 11215
<< metal4 >>
rect 72947 19632 74630 21315
use cap_200p  cap_200p_0
timestamp 1668357910
transform 1 0 44238 0 1 22632
box -3186 -3040 60524 67041
use r_8k  r_8k_1
timestamp 1668357910
transform 1 0 72736 0 1 8422
box -2962 -2369 2460 2830
<< labels >>
rlabel metal2 71224 10791 71794 11361 0 vfine
port 1 n
rlabel metal3 73440 12603 74458 13621 7 vout
port 2 n
rlabel metal4 72947 19632 74630 21315 0 vss
port 3 n
rlabel metal2 69774 6219 70206 6651 7 vss
<< end >>
