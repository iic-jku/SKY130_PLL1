magic
tech sky130A
magscale 1 2
timestamp 1668357910
<< nwell >>
rect -1319 -289 1319 289
<< pmos >>
rect -1119 -70 -1089 70
rect -1023 -70 -993 70
rect -927 -70 -897 70
rect -831 -70 -801 70
rect -735 -70 -705 70
rect -639 -70 -609 70
rect -543 -70 -513 70
rect -447 -70 -417 70
rect -351 -70 -321 70
rect -255 -70 -225 70
rect -159 -70 -129 70
rect -63 -70 -33 70
rect 33 -70 63 70
rect 129 -70 159 70
rect 225 -70 255 70
rect 321 -70 351 70
rect 417 -70 447 70
rect 513 -70 543 70
rect 609 -70 639 70
rect 705 -70 735 70
rect 801 -70 831 70
rect 897 -70 927 70
rect 993 -70 1023 70
rect 1089 -70 1119 70
<< pdiff >>
rect -1181 58 -1119 70
rect -1181 -58 -1169 58
rect -1135 -58 -1119 58
rect -1181 -70 -1119 -58
rect -1089 58 -1023 70
rect -1089 -58 -1073 58
rect -1039 -58 -1023 58
rect -1089 -70 -1023 -58
rect -993 58 -927 70
rect -993 -58 -977 58
rect -943 -58 -927 58
rect -993 -70 -927 -58
rect -897 58 -831 70
rect -897 -58 -881 58
rect -847 -58 -831 58
rect -897 -70 -831 -58
rect -801 58 -735 70
rect -801 -58 -785 58
rect -751 -58 -735 58
rect -801 -70 -735 -58
rect -705 58 -639 70
rect -705 -58 -689 58
rect -655 -58 -639 58
rect -705 -70 -639 -58
rect -609 58 -543 70
rect -609 -58 -593 58
rect -559 -58 -543 58
rect -609 -70 -543 -58
rect -513 58 -447 70
rect -513 -58 -497 58
rect -463 -58 -447 58
rect -513 -70 -447 -58
rect -417 58 -351 70
rect -417 -58 -401 58
rect -367 -58 -351 58
rect -417 -70 -351 -58
rect -321 58 -255 70
rect -321 -58 -305 58
rect -271 -58 -255 58
rect -321 -70 -255 -58
rect -225 58 -159 70
rect -225 -58 -209 58
rect -175 -58 -159 58
rect -225 -70 -159 -58
rect -129 58 -63 70
rect -129 -58 -113 58
rect -79 -58 -63 58
rect -129 -70 -63 -58
rect -33 58 33 70
rect -33 -58 -17 58
rect 17 -58 33 58
rect -33 -70 33 -58
rect 63 58 129 70
rect 63 -58 79 58
rect 113 -58 129 58
rect 63 -70 129 -58
rect 159 58 225 70
rect 159 -58 175 58
rect 209 -58 225 58
rect 159 -70 225 -58
rect 255 58 321 70
rect 255 -58 271 58
rect 305 -58 321 58
rect 255 -70 321 -58
rect 351 58 417 70
rect 351 -58 367 58
rect 401 -58 417 58
rect 351 -70 417 -58
rect 447 58 513 70
rect 447 -58 463 58
rect 497 -58 513 58
rect 447 -70 513 -58
rect 543 58 609 70
rect 543 -58 559 58
rect 593 -58 609 58
rect 543 -70 609 -58
rect 639 58 705 70
rect 639 -58 655 58
rect 689 -58 705 58
rect 639 -70 705 -58
rect 735 58 801 70
rect 735 -58 751 58
rect 785 -58 801 58
rect 735 -70 801 -58
rect 831 58 897 70
rect 831 -58 847 58
rect 881 -58 897 58
rect 831 -70 897 -58
rect 927 58 993 70
rect 927 -58 943 58
rect 977 -58 993 58
rect 927 -70 993 -58
rect 1023 58 1089 70
rect 1023 -58 1039 58
rect 1073 -58 1089 58
rect 1023 -70 1089 -58
rect 1119 58 1181 70
rect 1119 -58 1135 58
rect 1169 -58 1181 58
rect 1119 -70 1181 -58
<< pdiffc >>
rect -1169 -58 -1135 58
rect -1073 -58 -1039 58
rect -977 -58 -943 58
rect -881 -58 -847 58
rect -785 -58 -751 58
rect -689 -58 -655 58
rect -593 -58 -559 58
rect -497 -58 -463 58
rect -401 -58 -367 58
rect -305 -58 -271 58
rect -209 -58 -175 58
rect -113 -58 -79 58
rect -17 -58 17 58
rect 79 -58 113 58
rect 175 -58 209 58
rect 271 -58 305 58
rect 367 -58 401 58
rect 463 -58 497 58
rect 559 -58 593 58
rect 655 -58 689 58
rect 751 -58 785 58
rect 847 -58 881 58
rect 943 -58 977 58
rect 1039 -58 1073 58
rect 1135 -58 1169 58
<< nsubdiff >>
rect -1283 219 -1187 253
rect 1187 219 1283 253
rect -1283 157 -1249 219
rect 1249 157 1283 219
rect -1283 -219 -1249 -157
rect 1249 -219 1283 -157
rect -1283 -253 -1187 -219
rect 1187 -253 1283 -219
<< nsubdiffcont >>
rect -1187 219 1187 253
rect -1283 -157 -1249 157
rect 1249 -157 1283 157
rect -1187 -253 1187 -219
<< poly >>
rect -1137 151 -1071 167
rect -1137 117 -1121 151
rect -1087 117 -1071 151
rect -1137 101 -1071 117
rect 1071 151 1137 167
rect 1071 117 1087 151
rect 1121 117 1137 151
rect 1071 101 1137 117
rect -1119 70 -1089 101
rect -1023 70 -993 97
rect -927 70 -897 97
rect -831 70 -801 97
rect -735 70 -705 97
rect -639 70 -609 97
rect -543 70 -513 97
rect -447 70 -417 97
rect -351 70 -321 97
rect -255 70 -225 97
rect -159 70 -129 97
rect -63 70 -33 97
rect 33 70 63 97
rect 129 70 159 97
rect 225 70 255 97
rect 321 70 351 97
rect 417 70 447 97
rect 513 70 543 97
rect 609 70 639 97
rect 705 70 735 97
rect 801 70 831 97
rect 897 70 927 96
rect 993 70 1023 96
rect 1089 70 1119 101
rect -1119 -96 -1089 -70
rect -1023 -101 -993 -70
rect -927 -101 -897 -70
rect -831 -101 -801 -70
rect -735 -101 -705 -70
rect -639 -101 -609 -70
rect -543 -101 -513 -70
rect -447 -101 -417 -70
rect -351 -101 -321 -70
rect -255 -101 -225 -70
rect -159 -101 -129 -70
rect -63 -101 -33 -70
rect 33 -101 63 -70
rect 129 -101 159 -70
rect 225 -101 255 -70
rect 321 -101 351 -70
rect 417 -101 447 -70
rect 513 -101 543 -70
rect 609 -101 639 -70
rect 705 -101 735 -70
rect 801 -101 831 -70
rect 897 -101 927 -70
rect 993 -101 1023 -70
rect 1089 -97 1119 -70
rect -1041 -117 1041 -101
rect -1041 -151 -1025 -117
rect -991 -151 -929 -117
rect -895 -151 -833 -117
rect -799 -151 -737 -117
rect -703 -151 -641 -117
rect -607 -151 -545 -117
rect -511 -151 -449 -117
rect -415 -151 -353 -117
rect -319 -151 -257 -117
rect -223 -151 -161 -117
rect -127 -151 -65 -117
rect -31 -151 31 -117
rect 65 -151 127 -117
rect 161 -151 223 -117
rect 257 -151 319 -117
rect 353 -151 415 -117
rect 449 -151 511 -117
rect 545 -151 607 -117
rect 641 -151 703 -117
rect 737 -151 799 -117
rect 833 -151 895 -117
rect 929 -151 991 -117
rect 1025 -151 1041 -117
rect -1041 -167 1041 -151
<< polycont >>
rect -1121 117 -1087 151
rect 1087 117 1121 151
rect -1025 -151 -991 -117
rect -929 -151 -895 -117
rect -833 -151 -799 -117
rect -737 -151 -703 -117
rect -641 -151 -607 -117
rect -545 -151 -511 -117
rect -449 -151 -415 -117
rect -353 -151 -319 -117
rect -257 -151 -223 -117
rect -161 -151 -127 -117
rect -65 -151 -31 -117
rect 31 -151 65 -117
rect 127 -151 161 -117
rect 223 -151 257 -117
rect 319 -151 353 -117
rect 415 -151 449 -117
rect 511 -151 545 -117
rect 607 -151 641 -117
rect 703 -151 737 -117
rect 799 -151 833 -117
rect 895 -151 929 -117
rect 991 -151 1025 -117
<< locali >>
rect -1283 219 -1187 253
rect 1187 219 1283 253
rect -1283 157 -1249 219
rect -1169 151 -1135 219
rect 1135 151 1169 219
rect -1169 117 -1121 151
rect -1087 117 -1071 151
rect 1071 117 1087 151
rect 1121 117 1169 151
rect -1169 58 -1135 117
rect -1169 -74 -1135 -58
rect -1073 58 -1039 74
rect -1073 -74 -1039 -58
rect -977 58 -943 74
rect -977 -74 -943 -58
rect -881 58 -847 74
rect -881 -74 -847 -58
rect -785 58 -751 74
rect -785 -74 -751 -58
rect -689 58 -655 74
rect -689 -74 -655 -58
rect -593 58 -559 74
rect -593 -74 -559 -58
rect -497 58 -463 74
rect -497 -74 -463 -58
rect -401 58 -367 74
rect -401 -74 -367 -58
rect -305 58 -271 74
rect -305 -74 -271 -58
rect -209 58 -175 74
rect -209 -74 -175 -58
rect -113 58 -79 74
rect -113 -74 -79 -58
rect -17 58 17 74
rect -17 -74 17 -58
rect 79 58 113 74
rect 79 -74 113 -58
rect 175 58 209 74
rect 175 -74 209 -58
rect 271 58 305 74
rect 271 -74 305 -58
rect 367 58 401 74
rect 367 -74 401 -58
rect 463 58 497 74
rect 463 -74 497 -58
rect 559 58 593 74
rect 559 -74 593 -58
rect 655 58 689 74
rect 655 -74 689 -58
rect 751 58 785 74
rect 751 -74 785 -58
rect 847 58 881 74
rect 847 -74 881 -58
rect 943 58 977 74
rect 943 -74 977 -58
rect 1039 58 1073 74
rect 1039 -74 1073 -58
rect 1135 58 1169 117
rect 1135 -74 1169 -58
rect 1249 157 1283 219
rect -1283 -219 -1249 -157
rect -1041 -117 1041 -109
rect -1041 -151 -1025 -117
rect -991 -151 -929 -117
rect -895 -151 -833 -117
rect -799 -151 -737 -117
rect -703 -151 -641 -117
rect -607 -151 -545 -117
rect -511 -151 -449 -117
rect -415 -151 -353 -117
rect -319 -151 -257 -117
rect -223 -151 -161 -117
rect -127 -151 -65 -117
rect -31 -151 31 -117
rect 65 -151 127 -117
rect 161 -151 223 -117
rect 257 -151 319 -117
rect 353 -151 415 -117
rect 449 -151 511 -117
rect 545 -151 607 -117
rect 641 -151 703 -117
rect 737 -151 799 -117
rect 833 -151 895 -117
rect 929 -151 991 -117
rect 1025 -151 1041 -117
rect -1041 -159 1041 -151
rect 1249 -219 1283 -157
rect -1283 -253 -1187 -219
rect 1187 -253 1283 -219
<< viali >>
rect -1121 117 -1087 151
rect 1087 117 1121 151
rect -1169 -58 -1135 58
rect -1073 -58 -1039 58
rect -977 -58 -943 58
rect -881 -58 -847 58
rect -785 -58 -751 58
rect -689 -58 -655 58
rect -593 -58 -559 58
rect -497 -58 -463 58
rect -401 -58 -367 58
rect -305 -58 -271 58
rect -209 -58 -175 58
rect -113 -58 -79 58
rect -17 -58 17 58
rect 79 -58 113 58
rect 175 -58 209 58
rect 271 -58 305 58
rect 367 -58 401 58
rect 463 -58 497 58
rect 559 -58 593 58
rect 655 -58 689 58
rect 751 -58 785 58
rect 847 -58 881 58
rect 943 -58 977 58
rect 1039 -58 1073 58
rect 1135 -58 1169 58
rect -1025 -151 -991 -117
rect -929 -151 -895 -117
rect -833 -151 -799 -117
rect -737 -151 -703 -117
rect -641 -151 -607 -117
rect -545 -151 -511 -117
rect -449 -151 -415 -117
rect -353 -151 -319 -117
rect -257 -151 -223 -117
rect -161 -151 -127 -117
rect -65 -151 -31 -117
rect 31 -151 65 -117
rect 127 -151 161 -117
rect 223 -151 257 -117
rect 319 -151 353 -117
rect 415 -151 449 -117
rect 511 -151 545 -117
rect 607 -151 641 -117
rect 703 -151 737 -117
rect 799 -151 833 -117
rect 895 -151 929 -117
rect 991 -151 1025 -117
<< metal1 >>
rect -1169 151 -1075 157
rect -1169 117 -1121 151
rect -1087 117 -1075 151
rect -1169 111 -1075 117
rect 1075 151 1169 157
rect 1075 117 1087 151
rect 1121 117 1169 151
rect 1075 111 1169 117
rect -1169 70 -1133 111
rect 1133 70 1169 111
rect -1180 63 -1028 70
rect -1180 7 -1179 63
rect -1126 7 -1083 63
rect -1030 7 -1028 63
rect -1180 0 -1169 7
rect -1175 -58 -1169 0
rect -1135 0 -1073 7
rect -1135 -58 -1129 0
rect -1175 -70 -1129 -58
rect -1079 -58 -1073 0
rect -1039 0 -1028 7
rect -983 58 -937 70
rect -983 0 -977 58
rect -1039 -58 -1033 0
rect -1079 -70 -1033 -58
rect -988 -7 -977 0
rect -943 0 -937 58
rect -892 63 -836 70
rect -892 7 -891 63
rect -838 7 -836 63
rect -892 0 -881 7
rect -943 -7 -932 0
rect -988 -63 -987 -7
rect -934 -63 -932 -7
rect -988 -70 -932 -63
rect -887 -58 -881 0
rect -847 0 -836 7
rect -791 58 -745 70
rect -791 0 -785 58
rect -847 -58 -841 0
rect -887 -70 -841 -58
rect -796 -7 -785 0
rect -751 0 -745 58
rect -700 63 -644 70
rect -700 7 -699 63
rect -646 7 -644 63
rect -700 0 -689 7
rect -751 -7 -740 0
rect -796 -63 -795 -7
rect -742 -63 -740 -7
rect -796 -70 -740 -63
rect -695 -58 -689 0
rect -655 0 -644 7
rect -599 58 -553 70
rect -599 0 -593 58
rect -655 -58 -649 0
rect -695 -70 -649 -58
rect -604 -7 -593 0
rect -559 0 -553 58
rect -508 63 -452 70
rect -508 7 -507 63
rect -454 7 -452 63
rect -508 0 -497 7
rect -559 -7 -548 0
rect -604 -63 -603 -7
rect -550 -63 -548 -7
rect -604 -70 -548 -63
rect -503 -58 -497 0
rect -463 0 -452 7
rect -407 58 -361 70
rect -407 0 -401 58
rect -463 -58 -457 0
rect -503 -70 -457 -58
rect -412 -7 -401 0
rect -367 0 -361 58
rect -316 63 -260 70
rect -316 7 -315 63
rect -262 7 -260 63
rect -316 0 -305 7
rect -367 -7 -356 0
rect -412 -63 -411 -7
rect -358 -63 -356 -7
rect -412 -70 -356 -63
rect -311 -58 -305 0
rect -271 0 -260 7
rect -215 58 -169 70
rect -215 0 -209 58
rect -271 -58 -265 0
rect -311 -70 -265 -58
rect -220 -7 -209 0
rect -175 0 -169 58
rect -124 63 -68 70
rect -124 7 -123 63
rect -70 7 -68 63
rect -124 0 -113 7
rect -175 -7 -164 0
rect -220 -63 -219 -7
rect -166 -63 -164 -7
rect -220 -70 -164 -63
rect -119 -58 -113 0
rect -79 0 -68 7
rect -23 58 23 70
rect -23 0 -17 58
rect -79 -58 -73 0
rect -119 -70 -73 -58
rect -28 -7 -17 0
rect 17 0 23 58
rect 68 63 124 70
rect 68 7 69 63
rect 122 7 124 63
rect 68 0 79 7
rect 17 -7 28 0
rect -28 -63 -27 -7
rect 26 -63 28 -7
rect -28 -70 28 -63
rect 73 -58 79 0
rect 113 0 124 7
rect 169 58 215 70
rect 169 0 175 58
rect 113 -58 119 0
rect 73 -70 119 -58
rect 164 -7 175 0
rect 209 0 215 58
rect 260 63 316 70
rect 260 7 261 63
rect 314 7 316 63
rect 260 0 271 7
rect 209 -7 220 0
rect 164 -63 165 -7
rect 218 -63 220 -7
rect 164 -70 220 -63
rect 265 -58 271 0
rect 305 0 316 7
rect 361 58 407 70
rect 361 0 367 58
rect 305 -58 311 0
rect 265 -70 311 -58
rect 356 -7 367 0
rect 401 0 407 58
rect 452 63 508 70
rect 452 7 453 63
rect 506 7 508 63
rect 452 0 463 7
rect 401 -7 412 0
rect 356 -63 357 -7
rect 410 -63 412 -7
rect 356 -70 412 -63
rect 457 -58 463 0
rect 497 0 508 7
rect 553 58 599 70
rect 553 0 559 58
rect 497 -58 503 0
rect 457 -70 503 -58
rect 548 -7 559 0
rect 593 0 599 58
rect 644 63 700 70
rect 644 7 645 63
rect 698 7 700 63
rect 644 0 655 7
rect 593 -7 604 0
rect 548 -63 549 -7
rect 602 -63 604 -7
rect 548 -70 604 -63
rect 649 -58 655 0
rect 689 0 700 7
rect 745 58 791 70
rect 745 0 751 58
rect 689 -58 695 0
rect 649 -70 695 -58
rect 740 -7 751 0
rect 785 0 791 58
rect 836 63 892 70
rect 836 7 837 63
rect 890 7 892 63
rect 836 0 847 7
rect 785 -7 796 0
rect 740 -63 741 -7
rect 794 -63 796 -7
rect 740 -70 796 -63
rect 841 -58 847 0
rect 881 0 892 7
rect 937 58 983 70
rect 881 -58 887 0
rect 841 -70 887 -58
rect 937 -58 943 58
rect 977 -58 983 58
rect 1028 63 1180 70
rect 1028 7 1029 63
rect 1082 7 1125 63
rect 1178 7 1180 63
rect 1028 0 1039 7
rect 937 -109 983 -58
rect 1033 -58 1039 0
rect 1073 0 1135 7
rect 1073 -58 1079 0
rect 1033 -70 1079 -58
rect 1129 -58 1135 0
rect 1169 0 1180 7
rect 1169 -58 1175 0
rect 1129 -70 1175 -58
rect -1041 -117 1041 -109
rect -1041 -151 -1025 -117
rect -991 -151 -929 -117
rect -895 -151 -833 -117
rect -799 -151 -737 -117
rect -703 -151 -641 -117
rect -607 -151 -545 -117
rect -511 -151 -449 -117
rect -415 -151 -353 -117
rect -319 -151 -257 -117
rect -223 -151 -161 -117
rect -127 -151 -65 -117
rect -31 -151 31 -117
rect 65 -151 127 -117
rect 161 -151 223 -117
rect 257 -151 319 -117
rect 353 -151 415 -117
rect 449 -151 511 -117
rect 545 -151 607 -117
rect 641 -151 703 -117
rect 737 -151 799 -117
rect 833 -151 895 -117
rect 929 -151 991 -117
rect 1025 -151 1041 -117
rect -1041 -159 1041 -151
<< via1 >>
rect -1179 58 -1126 63
rect -1179 7 -1169 58
rect -1169 7 -1135 58
rect -1135 7 -1126 58
rect -1083 58 -1030 63
rect -1083 7 -1073 58
rect -1073 7 -1039 58
rect -1039 7 -1030 58
rect -891 58 -838 63
rect -891 7 -881 58
rect -881 7 -847 58
rect -847 7 -838 58
rect -987 -58 -977 -7
rect -977 -58 -943 -7
rect -943 -58 -934 -7
rect -987 -63 -934 -58
rect -699 58 -646 63
rect -699 7 -689 58
rect -689 7 -655 58
rect -655 7 -646 58
rect -795 -58 -785 -7
rect -785 -58 -751 -7
rect -751 -58 -742 -7
rect -795 -63 -742 -58
rect -507 58 -454 63
rect -507 7 -497 58
rect -497 7 -463 58
rect -463 7 -454 58
rect -603 -58 -593 -7
rect -593 -58 -559 -7
rect -559 -58 -550 -7
rect -603 -63 -550 -58
rect -315 58 -262 63
rect -315 7 -305 58
rect -305 7 -271 58
rect -271 7 -262 58
rect -411 -58 -401 -7
rect -401 -58 -367 -7
rect -367 -58 -358 -7
rect -411 -63 -358 -58
rect -123 58 -70 63
rect -123 7 -113 58
rect -113 7 -79 58
rect -79 7 -70 58
rect -219 -58 -209 -7
rect -209 -58 -175 -7
rect -175 -58 -166 -7
rect -219 -63 -166 -58
rect 69 58 122 63
rect 69 7 79 58
rect 79 7 113 58
rect 113 7 122 58
rect -27 -58 -17 -7
rect -17 -58 17 -7
rect 17 -58 26 -7
rect -27 -63 26 -58
rect 261 58 314 63
rect 261 7 271 58
rect 271 7 305 58
rect 305 7 314 58
rect 165 -58 175 -7
rect 175 -58 209 -7
rect 209 -58 218 -7
rect 165 -63 218 -58
rect 453 58 506 63
rect 453 7 463 58
rect 463 7 497 58
rect 497 7 506 58
rect 357 -58 367 -7
rect 367 -58 401 -7
rect 401 -58 410 -7
rect 357 -63 410 -58
rect 645 58 698 63
rect 645 7 655 58
rect 655 7 689 58
rect 689 7 698 58
rect 549 -58 559 -7
rect 559 -58 593 -7
rect 593 -58 602 -7
rect 549 -63 602 -58
rect 837 58 890 63
rect 837 7 847 58
rect 847 7 881 58
rect 881 7 890 58
rect 741 -58 751 -7
rect 751 -58 785 -7
rect 785 -58 794 -7
rect 741 -63 794 -58
rect 1029 58 1082 63
rect 1029 7 1039 58
rect 1039 7 1073 58
rect 1073 7 1082 58
rect 1125 58 1178 63
rect 1125 7 1135 58
rect 1135 7 1169 58
rect 1169 7 1178 58
<< metal2 >>
rect -1180 63 1180 70
rect -1180 7 -1179 63
rect -1126 7 -1083 63
rect -1030 28 -891 63
rect -1030 7 -1028 28
rect -1180 0 -1028 7
rect -892 7 -891 28
rect -838 28 -699 63
rect -838 7 -836 28
rect -892 0 -836 7
rect -700 7 -699 28
rect -646 28 -507 63
rect -646 7 -644 28
rect -700 0 -644 7
rect -508 7 -507 28
rect -454 28 -315 63
rect -454 7 -452 28
rect -508 0 -452 7
rect -316 7 -315 28
rect -262 28 -123 63
rect -262 7 -260 28
rect -316 0 -260 7
rect -124 7 -123 28
rect -70 28 69 63
rect -70 7 -68 28
rect -124 0 -68 7
rect 68 7 69 28
rect 122 28 261 63
rect 122 7 124 28
rect 68 0 124 7
rect 260 7 261 28
rect 314 28 453 63
rect 314 7 316 28
rect 260 0 316 7
rect 452 7 453 28
rect 506 28 645 63
rect 506 7 508 28
rect 452 0 508 7
rect 644 7 645 28
rect 698 28 837 63
rect 698 7 700 28
rect 644 0 700 7
rect 836 7 837 28
rect 890 28 1029 63
rect 890 7 892 28
rect 836 0 892 7
rect 1028 7 1029 28
rect 1082 7 1125 63
rect 1178 7 1180 63
rect 1028 0 1180 7
rect -988 -7 -932 0
rect -988 -28 -987 -7
rect -993 -63 -987 -28
rect -934 -28 -932 -7
rect -796 -7 -740 0
rect -796 -28 -795 -7
rect -934 -63 -795 -28
rect -742 -28 -740 -7
rect -604 -7 -548 0
rect -604 -28 -603 -7
rect -742 -63 -603 -28
rect -550 -28 -548 -7
rect -412 -7 -356 0
rect -412 -28 -411 -7
rect -550 -63 -411 -28
rect -358 -28 -356 -7
rect -220 -7 -164 0
rect -220 -28 -219 -7
rect -358 -63 -219 -28
rect -166 -28 -164 -7
rect -28 -7 28 0
rect -28 -28 -27 -7
rect -166 -63 -27 -28
rect 26 -28 28 -7
rect 164 -7 220 0
rect 164 -28 165 -7
rect 26 -63 165 -28
rect 218 -28 220 -7
rect 356 -7 412 0
rect 356 -28 357 -7
rect 218 -63 357 -28
rect 410 -28 412 -7
rect 548 -7 604 0
rect 548 -28 549 -7
rect 410 -63 549 -28
rect 602 -28 604 -7
rect 740 -7 796 0
rect 740 -28 741 -7
rect 602 -63 741 -28
rect 794 -28 796 -7
rect 794 -63 801 -28
rect -993 -70 801 -63
<< properties >>
string FIXED_BBOX -1266 -236 1266 236
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.7 l 0.15 m 1 nf 24 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
