magic
tech sky130A
magscale 1 2
timestamp 1669729258
<< metal1 >>
rect 26164 12562 26284 12568
rect -12163 12442 -5653 12562
rect -5533 12442 -5527 12562
rect 11722 12442 26164 12562
rect -12163 10339 -12043 12442
rect 26164 12436 26284 12442
rect -2464 10228 -2458 10528
rect -2158 10228 -2152 10528
rect 849 9938 855 10539
rect 1456 9938 1462 10539
rect 9045 9933 9051 10534
rect 9652 9933 9658 10534
rect 11562 10228 11568 10528
rect 11868 10228 11874 10528
rect -20724 9290 -20624 9301
rect -5611 9190 -5605 9290
rect -5505 9190 -5498 9290
rect -20724 8422 -20624 9190
rect 1616 9154 1628 9755
rect 2229 9154 2235 9755
rect 8298 9167 8305 9768
rect 8906 9167 8912 9768
rect 14915 9146 14955 9338
rect -19756 8915 -19750 8967
rect -19698 8962 -19692 8967
rect -19698 8920 -19353 8962
rect -19698 8915 -19692 8920
rect -17182 8742 -17176 8794
rect -17124 8742 -17118 8794
rect -14914 7601 -14908 7653
rect -14856 7601 -14850 7653
rect -20699 6598 -20647 6604
rect -20647 6551 -19311 6593
rect -20699 6540 -20647 6546
rect -16102 5460 -14168 5530
rect -14210 5335 -14168 5460
rect -2038 3494 -1972 4835
rect 1620 3725 1632 4326
rect 2233 3725 2239 4326
rect 8281 3735 8293 4336
rect 8894 3735 8900 4336
rect 12016 4118 12022 4170
rect 12074 4118 12080 4170
rect -2038 3422 -1972 3428
rect -14023 3103 -14017 3169
rect -13951 3103 -13294 3169
rect 872 2983 878 3584
rect 1479 2983 1485 3584
rect 9069 2951 9075 3552
rect 9676 2951 9682 3552
rect 12445 -393 12515 -387
rect 12445 -538 12515 -463
rect -32592 -573 -32022 -558
rect -32592 -1111 -32348 -573
rect -32256 -1111 -32022 -573
rect -32592 -1128 -32022 -1111
rect -18372 -573 -18252 -558
rect -18372 -1111 -18358 -573
rect -18266 -1111 -18252 -573
rect -18372 -1128 -18252 -1111
rect -1340 -573 -770 -558
rect -1340 -1111 -1096 -573
rect -1004 -1111 -770 -573
rect -1340 -1128 -770 -1111
rect 5117 -932 5417 -926
rect 5117 -1243 5417 -1237
rect 4771 -2504 5763 -2408
rect 5626 -3741 5678 -3735
rect 4851 -3747 4857 -3741
rect 4811 -3787 4857 -3747
rect 4851 -3793 4857 -3787
rect 4909 -3793 4915 -3741
rect 5678 -3787 5724 -3747
rect 5626 -3799 5678 -3793
rect 5117 -4387 5417 -4381
rect 5117 -4693 5417 -4687
rect 3723 -9970 3789 -9964
rect 5977 -9970 6043 -9964
rect 3717 -10036 3723 -9970
rect 3789 -10036 5977 -9970
rect 3723 -10042 3789 -10036
rect 5977 -10042 6043 -10036
rect -44044 -11174 -43474 -10604
rect -42408 -11174 -41838 -10604
rect -40772 -11174 -40202 -10604
rect -39136 -11174 -38566 -10604
rect -37500 -11174 -36930 -10604
rect -35864 -11174 -35294 -10604
rect -34228 -11174 -33658 -10604
rect -32592 -11174 -32022 -10604
rect -30054 -11174 -29484 -10604
rect -28418 -11174 -27848 -10604
rect -26782 -11174 -26212 -10604
rect -25146 -11174 -24576 -10604
rect -23510 -11174 -22940 -10604
rect -21874 -11174 -21304 -10604
rect -20238 -11174 -19668 -10604
rect -18602 -11174 -18032 -10604
rect -16064 -11174 -15494 -10604
rect -14428 -11174 -13858 -10604
rect -12792 -11174 -12222 -10604
rect -11156 -11174 -10586 -10604
rect -9520 -11174 -8950 -10604
rect -7884 -11174 -7314 -10604
rect -6248 -11174 -5678 -10604
rect -4612 -11174 -4042 -10604
rect -2976 -11174 -2406 -10604
rect -1340 -11174 -770 -10604
rect 12172 -11154 12742 -10584
rect 13808 -11154 14378 -10584
rect 15444 -11140 16014 -10584
rect 15443 -11154 16014 -11140
rect 17080 -11154 17650 -10584
rect 18716 -11135 19286 -10584
rect 18715 -11154 19286 -11135
rect 20352 -11136 20922 -10584
rect 20351 -11154 20922 -11136
rect 21988 -11154 22558 -10584
rect 23624 -11154 24194 -10584
rect -44044 -57797 -43944 -11174
rect -42407 -57507 -42307 -11174
rect -40772 -57217 -40672 -11174
rect -39135 -56927 -39035 -11174
rect -37500 -56637 -37400 -11174
rect -35864 -56347 -35764 -11174
rect -34227 -56057 -34127 -11174
rect -32591 -55767 -32491 -11174
rect -30054 -11288 -29954 -11174
rect -30054 -11399 -29954 -11388
rect -28417 -11299 -28317 -11174
rect -28417 -11405 -28317 -11399
rect -26782 -11299 -26682 -11174
rect -26782 -11405 -26682 -11399
rect -25145 -11299 -25045 -11174
rect -25145 -11405 -25045 -11399
rect -23510 -11299 -23410 -11174
rect -23510 -11405 -23410 -11399
rect -21874 -11299 -21774 -11174
rect -21874 -11405 -21774 -11399
rect -20237 -11299 -20137 -11174
rect -20237 -11405 -20137 -11399
rect -18601 -11299 -18501 -11174
rect -18601 -11405 -18501 -11399
rect -16065 -11678 -15965 -11174
rect -26420 -11778 -15965 -11678
rect -26420 -13641 -26320 -11778
rect -14428 -11968 -14328 -11174
rect -23476 -12068 -14328 -11968
rect -23476 -13602 -23376 -12068
rect -12793 -12258 -12693 -11174
rect -23476 -13708 -23376 -13702
rect -20540 -12358 -12693 -12258
rect -20540 -13634 -20440 -12358
rect -11156 -12548 -11056 -11174
rect -20540 -13740 -20440 -13734
rect -17587 -12648 -11056 -12548
rect -17587 -13644 -17487 -12648
rect -9521 -12838 -9421 -11174
rect -26420 -13747 -26320 -13741
rect -17587 -13750 -17487 -13744
rect -14651 -12938 -9421 -12838
rect -14651 -13650 -14551 -12938
rect -7885 -13128 -7785 -11174
rect -14651 -13756 -14551 -13750
rect -11704 -13228 -7785 -13128
rect -11704 -13650 -11604 -13228
rect -8762 -13628 -8662 -13622
rect -6248 -13628 -6148 -11174
rect -8662 -13728 -6148 -13628
rect -5817 -13631 -5717 -13625
rect -4612 -13631 -4512 -11174
rect -2976 -13508 -2876 -11174
rect -2976 -13514 -2773 -13508
rect -2976 -13614 -2873 -13514
rect -1340 -13511 -1240 -11174
rect 74 -13511 174 -13505
rect -1340 -13611 74 -13511
rect -2873 -13620 -2773 -13614
rect 74 -13617 174 -13611
rect -8762 -13734 -8662 -13728
rect -5717 -13731 -4512 -13631
rect -5817 -13737 -5717 -13731
rect -11704 -13756 -11604 -13750
rect 12171 -26970 12271 -11154
rect 12171 -27079 12177 -26970
rect 12265 -27079 12271 -26970
rect 12171 -27093 12271 -27079
rect 13808 -30642 13908 -11154
rect 13808 -30751 13814 -30642
rect 13902 -30751 13908 -30642
rect 13808 -30765 13908 -30751
rect 15443 -34314 15543 -11154
rect 15443 -34423 15449 -34314
rect 15537 -34423 15543 -34314
rect 15443 -34437 15543 -34423
rect 17080 -37986 17180 -11154
rect 17080 -38095 17086 -37986
rect 17174 -38095 17180 -37986
rect 17080 -38109 17180 -38095
rect 18715 -41658 18815 -11154
rect 18715 -41767 18721 -41658
rect 18809 -41767 18815 -41658
rect 18715 -41780 18815 -41767
rect 20351 -45330 20451 -11154
rect 20351 -45439 20357 -45330
rect 20445 -45439 20451 -45330
rect 20351 -45453 20451 -45439
rect 21988 -49002 22088 -11154
rect 21988 -49111 21994 -49002
rect 22082 -49111 22088 -49002
rect 21988 -49125 22088 -49111
rect 23624 -52674 23724 -11154
rect 25008 -16069 25128 -15594
rect 26242 -16069 26362 -15594
rect 25008 -16189 26362 -16069
rect 23624 -52783 23630 -52674
rect 23718 -52783 23724 -52674
rect 23624 -52797 23724 -52783
rect -26701 -55767 -26601 -55761
rect -32591 -55867 -26701 -55767
rect -26701 -55873 -26601 -55867
rect -23940 -56057 -23840 -56051
rect -34227 -56157 -23940 -56057
rect -23940 -56163 -23840 -56157
rect -21176 -56347 -21076 -56341
rect -35864 -56447 -21176 -56347
rect -21176 -56453 -21076 -56447
rect -18424 -56637 -18324 -56631
rect -37500 -56737 -18424 -56637
rect -18424 -56743 -18324 -56737
rect -15667 -56927 -15567 -56921
rect -39135 -57027 -15667 -56927
rect -15667 -57033 -15567 -57027
rect -12906 -57217 -12806 -57211
rect -40772 -57317 -12906 -57217
rect -12906 -57323 -12806 -57317
rect -10139 -57507 -10039 -57501
rect -42407 -57607 -10139 -57507
rect -10139 -57613 -10039 -57607
rect -7381 -57797 -7281 -57791
rect -44044 -57897 -7381 -57797
rect -7381 -57903 -7281 -57897
<< via1 >>
rect -5653 12442 -5533 12562
rect 26164 12442 26284 12562
rect -2458 10228 -2158 10528
rect 855 9938 1456 10539
rect 9051 9933 9652 10534
rect 11568 10228 11868 10528
rect -20724 9190 -20624 9290
rect -5605 9190 -5505 9290
rect 1628 9154 2229 9755
rect 8305 9167 8906 9768
rect -19750 8915 -19698 8967
rect -17176 8742 -17124 8794
rect -14908 7601 -14856 7653
rect -20699 6546 -20647 6598
rect 1632 3725 2233 4326
rect 8293 3735 8894 4336
rect 12022 4118 12074 4170
rect -2038 3428 -1972 3494
rect -14017 3103 -13951 3169
rect 878 2983 1479 3584
rect 9075 2951 9676 3552
rect 12445 -463 12515 -393
rect -32348 -1111 -32256 -573
rect -18358 -1111 -18266 -573
rect -1096 -1111 -1004 -573
rect 5117 -1237 5417 -932
rect 4857 -3793 4909 -3741
rect 5626 -3793 5678 -3741
rect 5117 -4687 5417 -4387
rect 3723 -10036 3789 -9970
rect 5977 -10036 6043 -9970
rect -30054 -11388 -29954 -11288
rect -28417 -11399 -28317 -11299
rect -26782 -11399 -26682 -11299
rect -25145 -11399 -25045 -11299
rect -23510 -11399 -23410 -11299
rect -21874 -11399 -21774 -11299
rect -20237 -11399 -20137 -11299
rect -18601 -11399 -18501 -11299
rect -26420 -13741 -26320 -13641
rect -23476 -13702 -23376 -13602
rect -20540 -13734 -20440 -13634
rect -17587 -13744 -17487 -13644
rect -14651 -13750 -14551 -13650
rect -11704 -13750 -11604 -13650
rect -8762 -13728 -8662 -13628
rect -2873 -13614 -2773 -13514
rect 74 -13611 174 -13511
rect -5817 -13731 -5717 -13631
rect 12177 -27079 12265 -26970
rect 13814 -30751 13902 -30642
rect 15449 -34423 15537 -34314
rect 17086 -38095 17174 -37986
rect 18721 -41767 18809 -41658
rect 20357 -45439 20445 -45330
rect 21994 -49111 22082 -49002
rect 23630 -52783 23718 -52674
rect -26701 -55867 -26601 -55767
rect -23940 -56157 -23840 -56057
rect -21176 -56447 -21076 -56347
rect -18424 -56737 -18324 -56637
rect -15667 -57027 -15567 -56927
rect -12906 -57317 -12806 -57217
rect -10139 -57607 -10039 -57507
rect -7381 -57897 -7281 -57797
<< metal2 >>
rect 9343 13130 9643 13139
rect 9643 12830 10136 12900
rect 9343 12821 9643 12830
rect -5653 12562 -5533 12568
rect -5533 12442 10661 12562
rect 26158 12442 26164 12562
rect 26284 12442 26290 12562
rect -5653 12436 -5533 12442
rect 9342 12261 9642 12270
rect 9333 11961 9342 12261
rect 9642 12191 10328 12261
rect 9642 11961 9651 12191
rect 9342 11952 9642 11961
rect -12681 10899 -12381 10908
rect -11821 10599 -11812 10899
rect -11512 10599 -11503 10899
rect -12681 10590 -12381 10599
rect -12451 10142 -12381 10590
rect -11812 10238 -11742 10599
rect 855 10539 1456 10545
rect -2458 10528 -2158 10534
rect -2467 10228 -2458 10528
rect -2158 10228 -2149 10528
rect -2458 10222 -2158 10228
rect -2467 9687 -2458 9987
rect -2158 9687 -2149 9987
rect 846 9938 855 10539
rect 1456 9938 1465 10539
rect 9051 10534 9652 10543
rect 855 9932 1456 9938
rect 11568 10528 11868 10534
rect 11559 10228 11568 10528
rect 11868 10228 11877 10528
rect 11568 10222 11868 10228
rect 9051 9924 9652 9933
rect 8305 9768 8906 9774
rect 1628 9755 2229 9761
rect -20724 9290 -20624 9301
rect -5605 9290 -5505 9296
rect -7513 9190 -7504 9290
rect -7404 9190 -5605 9290
rect -20724 9181 -20624 9190
rect -5605 9184 -5505 9190
rect 1619 9154 1628 9755
rect 2229 9154 2238 9755
rect 8296 9167 8305 9768
rect 8906 9167 8915 9768
rect 11559 9687 11568 9987
rect 11868 9687 11877 9987
rect 8305 9161 8906 9167
rect 1628 9148 2229 9154
rect -17718 9058 -17709 9124
rect -17643 9058 -17634 9124
rect -19750 8971 -19698 8973
rect -19763 8911 -19754 8971
rect -19694 8911 -19685 8971
rect -17709 8920 -17643 9058
rect -19750 8909 -19698 8911
rect -17176 8798 -17124 8800
rect -17189 8738 -17180 8798
rect -17120 8738 -17111 8798
rect -17176 8736 -17124 8738
rect -19715 8631 -19415 8640
rect -15155 8401 -15146 8701
rect -14846 8401 -14837 8701
rect 12146 8684 12155 8713
rect 12069 8642 12155 8684
rect 12146 8613 12155 8642
rect 12255 8613 12264 8713
rect -13588 8422 -13288 8431
rect -19715 8322 -19415 8331
rect -21698 8091 -21330 8125
rect -13588 8113 -13288 8122
rect -21698 7791 -21659 8091
rect -21359 7791 -21023 8091
rect -19586 7992 -19516 7998
rect -21698 7757 -21330 7791
rect -14908 7657 -14856 7659
rect -14921 7597 -14912 7657
rect -14852 7597 -14843 7657
rect -14908 7595 -14856 7597
rect -20694 6598 -20652 6736
rect -20705 6546 -20699 6598
rect -20647 6546 -20641 6598
rect -20384 6296 -20314 6832
rect -16001 6659 -15992 6959
rect -15692 6659 -15683 6959
rect -11205 6717 -11196 6845
rect -11068 6717 -11059 6845
rect -1335 6717 -1326 6845
rect -1198 6717 -1189 6845
rect -20624 5996 -20615 6296
rect -20315 5996 -20306 6296
rect -18733 5760 -18433 5769
rect -18733 5451 -18433 5460
rect -11196 4796 -11068 6717
rect 12146 6636 12155 6665
rect 12069 6594 12155 6636
rect 12146 6565 12155 6594
rect 12255 6565 12264 6665
rect 12146 4588 12155 4617
rect 12069 4546 12155 4588
rect 12146 4517 12155 4546
rect 12255 4517 12264 4617
rect 8293 4336 8894 4342
rect 1632 4326 2233 4332
rect -2584 4094 -2284 4103
rect -2584 3785 -2284 3794
rect -1715 4094 -1415 4103
rect -1715 3785 -1415 3794
rect 1623 3725 1632 4326
rect 2233 3725 2242 4326
rect 8284 3735 8293 4336
rect 8894 3735 8903 4336
rect 12445 4179 12515 4188
rect 12013 4174 12445 4179
rect 12009 4170 12445 4174
rect 12009 4118 12022 4170
rect 12074 4118 12445 4170
rect 12009 4114 12445 4118
rect 12013 4109 12445 4114
rect 12445 4100 12515 4109
rect 8293 3729 8894 3735
rect 1632 3719 2233 3725
rect 878 3584 1479 3593
rect -2038 3494 -1972 3503
rect -2044 3428 -2038 3494
rect -1972 3428 -1966 3494
rect -2038 3419 -1972 3428
rect -29397 3376 -29297 3385
rect -20031 3376 -19931 3385
rect -29297 3276 -20031 3376
rect -14378 3298 -14369 3364
rect -14303 3298 -14088 3364
rect -29397 3267 -29297 3276
rect -20031 3267 -19931 3276
rect -28997 2976 -28897 2985
rect -19890 2976 -19790 2985
rect -28897 2876 -19890 2976
rect -15372 2903 -15363 3203
rect -15063 2903 -15054 3203
rect -14154 3169 -14088 3298
rect -11800 3340 -11500 3349
rect -14017 3169 -13951 3175
rect -14154 3103 -14017 3169
rect -14017 3097 -13951 3103
rect -11800 3031 -11500 3040
rect 878 2974 1479 2983
rect 9075 3552 9676 3561
rect 9075 2942 9676 2951
rect -28997 2867 -28897 2876
rect -19890 2867 -19790 2876
rect 11099 2655 11169 3331
rect 10869 2646 11169 2655
rect 11738 2646 11808 3240
rect -28597 2576 -28497 2585
rect -19749 2576 -19649 2585
rect -28497 2476 -19749 2576
rect -28597 2467 -28497 2476
rect -19749 2467 -19649 2476
rect 11729 2346 11738 2646
rect 12038 2346 12047 2646
rect 10869 2337 11169 2346
rect -16842 2298 -16542 2307
rect -16542 1998 -16084 2068
rect -16842 1989 -16542 1998
rect -2869 1707 -2860 2139
rect -2428 1707 -2419 2139
rect 12445 1730 12515 1739
rect 12445 -393 12515 1660
rect 12439 -463 12445 -393
rect 12515 -463 12521 -393
rect 12445 -472 12515 -463
rect -32362 -573 -32242 -558
rect -32362 -1111 -32348 -573
rect -32256 -1111 -32242 -573
rect -32362 -1128 -32242 -1111
rect -18372 -573 -18252 -558
rect -18372 -1111 -18358 -573
rect -18266 -1111 -18252 -573
rect -18372 -1128 -18252 -1111
rect -1110 -573 -990 -558
rect -1110 -1111 -1096 -573
rect -1004 -1111 -990 -573
rect 5117 -932 5417 -923
rect -1110 -1128 -990 -1111
rect 5111 -1237 5117 -932
rect 5417 -1237 5423 -932
rect 5117 -1246 5417 -1237
rect 4853 -3737 4913 -3728
rect 5622 -3737 5682 -3728
rect 5620 -3793 5622 -3741
rect 5682 -3793 5684 -3741
rect 4853 -3806 4913 -3797
rect 5622 -3806 5682 -3797
rect 5117 -4387 5417 -4378
rect 5111 -4687 5117 -4387
rect 5417 -4687 5423 -4387
rect 5117 -4696 5417 -4687
rect -45469 -6464 -45460 -6032
rect -45028 -6464 -45019 -6032
rect 25169 -6444 25178 -6012
rect 25610 -6444 25619 -6012
rect 3723 -9970 3789 -9964
rect 3714 -10036 3723 -9970
rect 3789 -10036 3798 -9970
rect 5971 -10036 5977 -9970
rect 6043 -10036 6049 -9970
rect 3723 -10042 3789 -10036
rect -30060 -11388 -30054 -11288
rect -29954 -11388 -29948 -11288
rect -32018 -11488 -29954 -11388
rect -28423 -11399 -28417 -11299
rect -28317 -11399 -28311 -11299
rect -26788 -11399 -26782 -11299
rect -26682 -11399 -26676 -11299
rect -25151 -11399 -25145 -11299
rect -25045 -11399 -25039 -11299
rect -23516 -11399 -23510 -11299
rect -23410 -11399 -23404 -11299
rect -21880 -11399 -21874 -11299
rect -21774 -11399 -21768 -11299
rect -20243 -11399 -20237 -11299
rect -20137 -11399 -20131 -11299
rect -18607 -11399 -18601 -11299
rect -18501 -11399 -18495 -11299
rect -32018 -52673 -31918 -11488
rect -28417 -11678 -28317 -11399
rect -31728 -11778 -28317 -11678
rect -31728 -49001 -31628 -11778
rect -26782 -11968 -26682 -11399
rect -31438 -12068 -26682 -11968
rect -31438 -45329 -31338 -12068
rect -25145 -12258 -25045 -11399
rect -31148 -12358 -25045 -12258
rect -31148 -41657 -31048 -12358
rect -23510 -12548 -23410 -11399
rect -30858 -12648 -23410 -12548
rect -30858 -37985 -30758 -12648
rect -21874 -12838 -21774 -11399
rect -30568 -12938 -21774 -12838
rect -30568 -34313 -30468 -12938
rect -20237 -13128 -20137 -11399
rect -30278 -13228 -20137 -13128
rect -30278 -30641 -30178 -13228
rect -18601 -13418 -18501 -11399
rect -29988 -13518 -18501 -13418
rect -29988 -26969 -29888 -13518
rect -26426 -13741 -26420 -13641
rect -26320 -13741 -26314 -13641
rect -23482 -13702 -23476 -13602
rect -23376 -13702 -23370 -13602
rect -2879 -13614 -2873 -13514
rect -2773 -13614 -2767 -13514
rect 68 -13611 74 -13511
rect 174 -13611 180 -13511
rect 3027 -13584 3036 -13524
rect 3096 -13584 3105 -13524
rect -26402 -13889 -26346 -13741
rect -23458 -13863 -23402 -13702
rect -20546 -13734 -20540 -13634
rect -20440 -13734 -20434 -13634
rect -20514 -13889 -20458 -13734
rect -17593 -13744 -17587 -13644
rect -17487 -13744 -17481 -13644
rect -17570 -13863 -17514 -13744
rect -14657 -13750 -14651 -13650
rect -14551 -13750 -14545 -13650
rect -11710 -13750 -11704 -13650
rect -11604 -13750 -11598 -13650
rect -8768 -13728 -8762 -13628
rect -8662 -13728 -8656 -13628
rect -14626 -13863 -14570 -13750
rect -11682 -13863 -11626 -13750
rect -8738 -13871 -8682 -13728
rect -5823 -13731 -5817 -13631
rect -5717 -13731 -5711 -13631
rect -5794 -13863 -5738 -13731
rect -2850 -13863 -2794 -13614
rect 94 -13863 150 -13611
rect 3038 -13871 3094 -13584
rect 5977 -13867 6043 -10036
rect 25536 -12795 25836 -12786
rect 8900 -13600 25128 -13500
rect 8926 -13863 8982 -13600
rect 25008 -14534 25128 -13600
rect 25536 -13935 25836 -13095
rect 25396 -14005 25974 -13935
rect 26164 -14534 26284 12442
rect 24757 -16754 24827 -15834
rect 26543 -16754 26613 -15834
rect 24518 -17054 24527 -16754
rect 24827 -17054 24836 -16754
rect 26534 -17054 26543 -16754
rect 26843 -17054 26852 -16754
rect 12171 -26964 12271 -26955
rect -29988 -27079 -29984 -26969
rect -29892 -27079 -29888 -26969
rect -29988 -27094 -29888 -27079
rect 12162 -26970 12279 -26964
rect 12162 -27079 12177 -26970
rect 12265 -27079 12279 -26970
rect 12162 -27084 12279 -27079
rect 12171 -27093 12271 -27084
rect 13808 -30636 13908 -30627
rect -30278 -30751 -30274 -30641
rect -30182 -30751 -30178 -30641
rect -30278 -30766 -30178 -30751
rect 13799 -30642 13916 -30636
rect 13799 -30751 13814 -30642
rect 13902 -30751 13916 -30642
rect 13799 -30756 13916 -30751
rect 13808 -30765 13908 -30756
rect 15443 -34308 15543 -34299
rect -30568 -34423 -30564 -34313
rect -30472 -34423 -30468 -34313
rect -30568 -34438 -30468 -34423
rect 15434 -34314 15551 -34308
rect 15434 -34423 15449 -34314
rect 15537 -34423 15551 -34314
rect 15434 -34428 15551 -34423
rect 15443 -34437 15543 -34428
rect 17080 -37980 17180 -37971
rect -30858 -38095 -30854 -37985
rect -30762 -38095 -30758 -37985
rect -30858 -38110 -30758 -38095
rect 17071 -37986 17188 -37980
rect 17071 -38095 17086 -37986
rect 17174 -38095 17188 -37986
rect 17071 -38100 17188 -38095
rect 17080 -38109 17180 -38100
rect 18715 -41652 18815 -41643
rect -31148 -41767 -31144 -41657
rect -31052 -41767 -31048 -41657
rect -31148 -41782 -31048 -41767
rect 18706 -41658 18823 -41652
rect 18706 -41767 18721 -41658
rect 18809 -41767 18823 -41658
rect 18706 -41772 18823 -41767
rect 18715 -41781 18815 -41772
rect 20351 -45324 20451 -45315
rect -31438 -45439 -31434 -45329
rect -31342 -45439 -31338 -45329
rect -31438 -45454 -31338 -45439
rect 20342 -45330 20459 -45324
rect 20342 -45439 20357 -45330
rect 20445 -45439 20459 -45330
rect 20342 -45444 20459 -45439
rect 20351 -45453 20451 -45444
rect 21988 -48996 22088 -48987
rect -31728 -49111 -31724 -49001
rect -31632 -49111 -31628 -49001
rect -31728 -49126 -31628 -49111
rect 21979 -49002 22096 -48996
rect 21979 -49111 21994 -49002
rect 22082 -49111 22096 -49002
rect 21979 -49116 22096 -49111
rect 21988 -49125 22088 -49116
rect 23624 -52668 23724 -52659
rect -32018 -52783 -32014 -52673
rect -31922 -52783 -31918 -52673
rect -32018 -52798 -31918 -52783
rect 23615 -52674 23732 -52668
rect 23615 -52783 23630 -52674
rect 23718 -52783 23732 -52674
rect 23615 -52788 23732 -52783
rect 23624 -52797 23724 -52788
rect -26678 -54643 -26622 -54616
rect -28076 -54700 -26622 -54643
rect -26678 -54901 -26622 -54700
rect -23918 -54901 -23862 -54628
rect -21158 -54898 -21102 -54640
rect -18398 -54895 -18342 -54640
rect -26701 -55767 -26601 -54901
rect -26707 -55867 -26701 -55767
rect -26601 -55867 -26595 -55767
rect -23940 -56057 -23840 -54901
rect -23946 -56157 -23940 -56057
rect -23840 -56157 -23834 -56057
rect -21176 -56347 -21076 -54898
rect -21182 -56447 -21176 -56347
rect -21076 -56447 -21070 -56347
rect -18424 -56637 -18324 -54895
rect -15638 -54898 -15582 -54628
rect -12878 -54898 -12822 -54593
rect -18430 -56737 -18424 -56637
rect -18324 -56737 -18318 -56637
rect -15667 -56927 -15567 -54898
rect -15673 -57027 -15667 -56927
rect -15567 -57027 -15561 -56927
rect -12906 -57217 -12806 -54898
rect -10118 -54901 -10062 -54616
rect -7358 -54898 -7302 -54605
rect -4598 -54892 -4542 -54605
rect -1838 -54891 -1782 -54628
rect 922 -54890 978 -54628
rect -12912 -57317 -12906 -57217
rect -12806 -57317 -12800 -57217
rect -10139 -57507 -10039 -54901
rect -10145 -57607 -10139 -57507
rect -10039 -57607 -10033 -57507
rect -7381 -57797 -7281 -54898
rect -4622 -54901 -4522 -54892
rect -4622 -55010 -4522 -55001
rect -1860 -54900 -1760 -54891
rect -1860 -55009 -1760 -55000
rect 899 -54899 999 -54890
rect 3682 -54891 3738 -54628
rect 6442 -54891 6498 -54628
rect 9202 -54891 9258 -54628
rect 899 -55008 999 -54999
rect 3659 -54900 3759 -54891
rect 3659 -55009 3759 -55000
rect 6419 -54900 6519 -54891
rect 6419 -55009 6519 -55000
rect 9179 -54900 9279 -54891
rect 9179 -55009 9279 -55000
rect -7387 -57897 -7381 -57797
rect -7281 -57897 -7275 -57797
<< via2 >>
rect 9343 12830 9643 13130
rect 9342 11961 9642 12261
rect -12681 10599 -12381 10899
rect -11812 10599 -11512 10899
rect -2458 10228 -2158 10528
rect -2458 9687 -2158 9987
rect 855 9938 1456 10539
rect 9051 9933 9652 10534
rect 11568 10228 11868 10528
rect -20719 9195 -20629 9285
rect -7504 9190 -7404 9290
rect 1628 9154 2229 9755
rect 8305 9167 8906 9768
rect 11568 9687 11868 9987
rect -17709 9058 -17643 9124
rect -19754 8967 -19694 8971
rect -19754 8915 -19750 8967
rect -19750 8915 -19698 8967
rect -19698 8915 -19694 8967
rect -19754 8911 -19694 8915
rect -17180 8794 -17120 8798
rect -17180 8742 -17176 8794
rect -17176 8742 -17124 8794
rect -17124 8742 -17120 8794
rect -17180 8738 -17120 8742
rect -19715 8331 -19415 8631
rect -15146 8401 -14846 8701
rect 12155 8613 12255 8713
rect -13588 8122 -13288 8422
rect -21659 7791 -21359 8091
rect -14912 7653 -14852 7657
rect -14912 7601 -14908 7653
rect -14908 7601 -14856 7653
rect -14856 7601 -14852 7653
rect -14912 7597 -14852 7601
rect -15992 6659 -15692 6959
rect -11196 6717 -11068 6845
rect -1326 6717 -1198 6845
rect -20615 5996 -20315 6296
rect -18733 5460 -18433 5760
rect 12155 6565 12255 6665
rect -4426 6372 -3907 6499
rect 12155 4517 12255 4617
rect -2584 3794 -2284 4094
rect -1715 3794 -1415 4094
rect 1632 3725 2233 4326
rect 8293 3735 8894 4336
rect 12445 4109 12515 4179
rect -2038 3428 -1972 3494
rect -29397 3276 -29297 3376
rect -20031 3276 -19931 3376
rect -14369 3298 -14303 3364
rect -28997 2876 -28897 2976
rect -19890 2876 -19790 2976
rect -15363 2903 -15063 3203
rect -11800 3040 -11500 3340
rect 878 2983 1479 3584
rect 9075 2951 9676 3552
rect -28597 2476 -28497 2576
rect -19749 2476 -19649 2576
rect 10869 2346 11169 2646
rect 11738 2346 12038 2646
rect -16842 1998 -16542 2298
rect -2860 1707 -2428 2139
rect 12445 1660 12515 1730
rect -32348 -1111 -32256 -573
rect -18358 -1111 -18266 -573
rect -1096 -1111 -1004 -573
rect 5117 -1237 5417 -932
rect 4853 -3741 4913 -3737
rect 5622 -3741 5682 -3737
rect 4853 -3793 4857 -3741
rect 4857 -3793 4909 -3741
rect 4909 -3793 4913 -3741
rect 5622 -3793 5626 -3741
rect 5626 -3793 5678 -3741
rect 5678 -3793 5682 -3741
rect 4853 -3797 4913 -3793
rect 5622 -3797 5682 -3793
rect 5117 -4687 5417 -4387
rect -45460 -6464 -45028 -6032
rect 25178 -6444 25610 -6012
rect 3723 -10036 3789 -9970
rect 3036 -13584 3096 -13524
rect 25536 -13095 25836 -12795
rect 24527 -17054 24827 -16754
rect 26543 -17054 26843 -16754
rect -29984 -27079 -29892 -26969
rect 12177 -27079 12265 -26970
rect -30274 -30751 -30182 -30641
rect 13814 -30751 13902 -30642
rect -30564 -34423 -30472 -34313
rect 15449 -34423 15537 -34314
rect -30854 -38095 -30762 -37985
rect 17086 -38095 17174 -37986
rect -31144 -41767 -31052 -41657
rect 18721 -41767 18809 -41658
rect -31434 -45439 -31342 -45329
rect 20357 -45439 20445 -45330
rect -31724 -49111 -31632 -49001
rect 21994 -49111 22082 -49002
rect -32014 -52783 -31922 -52673
rect 23630 -52783 23718 -52674
rect -4622 -55001 -4522 -54901
rect -1860 -55000 -1760 -54900
rect 899 -54999 999 -54899
rect 3659 -55000 3759 -54900
rect 6419 -55000 6519 -54900
rect 9179 -55000 9279 -54900
<< metal3 >>
rect 9338 13135 9648 13141
rect 9338 12830 9343 12835
rect 9643 12830 9648 12835
rect 9338 12825 9648 12830
rect 9324 12261 9658 12277
rect 9324 11961 9342 12261
rect 9642 11961 9658 12261
rect 9324 11944 9658 11961
rect -12715 10899 -12347 10938
rect -12715 10599 -12681 10899
rect -12381 10599 -12347 10899
rect -12715 10570 -12347 10599
rect -11817 10899 -11807 10904
rect -11817 10599 -11812 10899
rect -11817 10594 -11807 10599
rect -11507 10594 -11501 10904
rect -2463 10528 -2453 10533
rect -2463 10228 -2458 10528
rect -2463 10223 -2453 10228
rect -2153 10223 -2147 10533
rect -2487 9987 -2119 10021
rect -2487 9687 -2458 9987
rect -2158 9687 -2119 9987
rect 844 9933 850 10544
rect 1451 10539 1461 10544
rect 1456 9938 1461 10539
rect 1451 9933 1461 9938
rect 9046 10534 9056 10539
rect 9046 9933 9051 10534
rect 9046 9928 9056 9933
rect 9657 9928 9663 10539
rect 11557 10223 11563 10533
rect 11863 10528 11873 10533
rect 11868 10228 11873 10528
rect 11863 10223 11873 10228
rect 11529 9987 11897 10021
rect -2487 9653 -2119 9687
rect 1623 9755 1633 9760
rect -20724 9290 -20624 9296
rect -7509 9290 -7399 9295
rect -20729 9285 -7504 9290
rect -20729 9195 -20719 9285
rect -20629 9195 -7504 9285
rect -20729 9190 -7504 9195
rect -7404 9190 -7399 9290
rect -20724 9185 -20624 9190
rect -7509 9185 -7399 9190
rect 1623 9154 1628 9755
rect 1623 9149 1633 9154
rect 2234 9149 2240 9760
rect 8294 9162 8300 9773
rect 8901 9768 8911 9773
rect 8906 9167 8911 9768
rect 11529 9687 11568 9987
rect 11868 9687 11897 9987
rect 11529 9653 11897 9687
rect 8901 9162 8911 9167
rect -17714 9124 -17638 9129
rect -32333 9058 -17709 9124
rect -17643 9058 -17638 9124
rect -32333 -558 -32267 9058
rect -17714 9053 -17638 9058
rect -19759 8971 -19689 8976
rect -19991 8911 -19754 8971
rect -19694 8911 -19689 8971
rect -21698 8091 -21330 8125
rect -21698 7791 -21659 8091
rect -21359 7791 -21330 8091
rect -21698 7757 -21330 7791
rect -20626 5991 -20620 6301
rect -20320 6296 -20310 6301
rect -20315 5996 -20310 6296
rect -20320 5991 -20310 5996
rect -19991 3381 -19931 8911
rect -19759 8906 -19689 8911
rect -17185 8798 -17115 8803
rect -19850 8738 -17180 8798
rect -17120 8738 -17115 8798
rect -29402 3376 -29292 3381
rect -29402 3276 -29397 3376
rect -29297 3276 -29292 3376
rect -29402 3271 -29292 3276
rect -20036 3376 -19926 3381
rect -20036 3276 -20031 3376
rect -19931 3276 -19926 3376
rect -20036 3271 -19926 3276
rect -32362 -573 -32242 -558
rect -32362 -1111 -32348 -573
rect -32256 -1111 -32242 -573
rect -32362 -1128 -32242 -1111
rect -45490 -6032 -45010 -6002
rect -45490 -6464 -45460 -6032
rect -45028 -6464 -45010 -6032
rect -45490 -6494 -45010 -6464
rect -29397 -23292 -29297 3271
rect -19850 2981 -19790 8738
rect -17185 8733 -17115 8738
rect 12150 8713 12260 8718
rect -15151 8701 -15141 8706
rect -19720 8631 -19410 8636
rect -19720 8626 -19715 8631
rect -19415 8626 -19410 8631
rect -15151 8401 -15146 8701
rect -15151 8396 -15141 8401
rect -14841 8396 -14835 8706
rect 12150 8613 12155 8713
rect 12255 8613 13715 8713
rect 12150 8608 12260 8613
rect -13622 8422 -13254 8461
rect -19720 8320 -19410 8326
rect -13622 8122 -13588 8422
rect -13288 8122 -13254 8422
rect -13622 8093 -13254 8122
rect -14917 7657 -14847 7662
rect -19709 7597 -14912 7657
rect -14852 7597 -14847 7657
rect -6094 7603 -105 7731
rect -29002 2976 -28892 2981
rect -29002 2876 -28997 2976
rect -28897 2876 -28892 2976
rect -29002 2871 -28892 2876
rect -19895 2976 -19785 2981
rect -19895 2876 -19890 2976
rect -19790 2876 -19785 2976
rect -19895 2871 -19785 2876
rect -28997 -19620 -28897 2871
rect -19709 2581 -19649 7597
rect -14917 7592 -14847 7597
rect -16021 6959 -15653 6993
rect -16021 6659 -15992 6959
rect -15692 6659 -15653 6959
rect -11201 6845 -11063 6850
rect -1331 6845 -1193 6850
rect -11201 6717 -11196 6845
rect -11068 6717 -1326 6845
rect -1198 6717 -1193 6845
rect -11201 6712 -11063 6717
rect -1331 6712 -1193 6717
rect -233 6715 -105 7603
rect -16021 6625 -15653 6659
rect 12150 6665 12260 6670
rect 12150 6565 12155 6665
rect 12255 6565 13315 6665
rect 12150 6560 12260 6565
rect -4449 6499 -3879 6525
rect -4449 6372 -4426 6499
rect -3907 6372 -3879 6499
rect -4449 6350 -3879 6372
rect -18767 5760 -18399 5789
rect -18767 5460 -18733 5760
rect -18433 5460 -18399 5760
rect -18767 5421 -18399 5460
rect -14374 3364 -14298 3369
rect -18343 3298 -14369 3364
rect -14303 3298 -14298 3364
rect -28602 2576 -28492 2581
rect -28602 2476 -28597 2576
rect -28497 2476 -28492 2576
rect -28602 2471 -28492 2476
rect -19754 2576 -19644 2581
rect -19754 2476 -19749 2576
rect -19649 2476 -19644 2576
rect -19754 2471 -19644 2476
rect -28597 -15948 -28497 2471
rect -18343 -558 -18277 3298
rect -14374 3293 -14298 3298
rect -11805 3345 -11495 3351
rect -15402 3203 -15034 3237
rect -15402 2903 -15363 3203
rect -15063 2903 -15034 3203
rect -11805 3040 -11800 3045
rect -11500 3040 -11495 3045
rect -11805 3035 -11495 3040
rect -15402 2869 -15034 2903
rect -16847 2303 -16537 2309
rect -16847 1998 -16842 2003
rect -16542 1998 -16537 2003
rect -16847 1993 -16537 1998
rect -4217 1304 -4151 6350
rect 12150 4617 12260 4622
rect 12150 4517 12155 4617
rect 12255 4517 12915 4617
rect 12150 4512 12260 4517
rect 8288 4336 8298 4341
rect 1627 4326 1637 4331
rect -2589 4094 -2279 4099
rect -2589 4089 -2584 4094
rect -2284 4089 -2279 4094
rect -2589 3783 -2279 3789
rect -1720 4094 -1410 4099
rect -1720 4089 -1715 4094
rect -1415 4089 -1410 4094
rect -1720 3783 -1410 3789
rect 1627 3725 1632 4326
rect 1627 3720 1637 3725
rect 2238 3720 2244 4331
rect 8288 3735 8293 4336
rect 8288 3730 8298 3735
rect 8899 3730 8905 4341
rect 12440 4179 12520 4184
rect 12440 4109 12445 4179
rect 12515 4109 12520 4179
rect 12440 4104 12520 4109
rect 873 3584 883 3589
rect -2043 3494 -1967 3499
rect -2043 3428 -2038 3494
rect -1972 3428 -1967 3494
rect -2043 3423 -1967 3428
rect -2038 2381 -1972 3423
rect 873 2983 878 3584
rect 873 2978 883 2983
rect 1484 2978 1490 3589
rect 9070 3552 9080 3557
rect 9070 2951 9075 3552
rect 9070 2946 9080 2951
rect 9681 2946 9687 3557
rect 10835 2646 11203 2675
rect -2038 2315 748 2381
rect -2865 2139 -2855 2144
rect -2865 1707 -2860 2139
rect -2865 1702 -2855 1707
rect -2423 1702 -2417 2144
rect -4217 1238 -1015 1304
rect -1081 -558 -1015 1238
rect -18372 -573 -18252 -558
rect -18372 -1111 -18358 -573
rect -18266 -1111 -18252 -573
rect -18372 -1128 -18252 -1111
rect -1110 -573 -990 -558
rect -1110 -1111 -1096 -573
rect -1004 -1111 -990 -573
rect -1110 -1128 -990 -1111
rect 682 -9970 748 2315
rect 10835 2346 10869 2646
rect 11169 2346 11203 2646
rect 10835 2307 11203 2346
rect 11733 2646 12043 2651
rect 11733 2641 11738 2646
rect 12038 2641 12043 2646
rect 11733 2335 12043 2341
rect 12445 1735 12515 4104
rect 12440 1730 12520 1735
rect 12440 1660 12445 1730
rect 12515 1660 12520 1730
rect 12440 1655 12520 1660
rect 5112 -927 5422 -921
rect 5112 -1237 5117 -1227
rect 5417 -1237 5422 -1227
rect 5112 -1242 5422 -1237
rect 4848 -3737 4918 -3732
rect 4848 -3797 4853 -3737
rect 4913 -3797 4918 -3737
rect 4848 -3802 4918 -3797
rect 5617 -3737 5687 -3732
rect 5617 -3797 5622 -3737
rect 5682 -3797 5687 -3737
rect 5617 -3802 5687 -3797
rect 3718 -9970 3794 -9965
rect 682 -10036 3723 -9970
rect 3789 -10036 3794 -9970
rect 3718 -10041 3794 -10036
rect 3031 -13524 3101 -13519
rect 4853 -13524 4913 -3802
rect 5083 -4387 5451 -4358
rect 5083 -4687 5117 -4387
rect 5417 -4687 5451 -4387
rect 5083 -4726 5451 -4687
rect 5622 -8680 5682 -3802
rect 3031 -13584 3036 -13524
rect 3096 -13584 4913 -13524
rect 3031 -13589 3101 -13584
rect 12815 -15948 12915 4517
rect -28597 -16068 -27956 -15948
rect 10553 -16068 12915 -15948
rect 13215 -19620 13315 6565
rect -28997 -19740 -27956 -19620
rect 10553 -19740 13315 -19620
rect 13615 -23292 13715 8613
rect 25151 -6012 25640 -5982
rect 25151 -6444 25178 -6012
rect 25610 -6444 25640 -6012
rect 25151 -6474 25640 -6444
rect 25531 -12790 25841 -12784
rect 25531 -13095 25536 -13090
rect 25836 -13095 25841 -13090
rect 25531 -13100 25841 -13095
rect 24498 -16754 24866 -16720
rect 24498 -17054 24527 -16754
rect 24827 -17054 24866 -16754
rect 24498 -17088 24866 -17054
rect 26504 -16754 26872 -16720
rect 26504 -17054 26543 -16754
rect 26843 -17054 26872 -16754
rect 26504 -17088 26872 -17054
rect -29397 -23412 -27956 -23292
rect 10506 -23412 13715 -23292
rect -29998 -26969 -27956 -26964
rect -29998 -27079 -29984 -26969
rect -29892 -27079 -27956 -26969
rect -29998 -27084 -27956 -27079
rect 10553 -26970 12286 -26964
rect 10553 -27079 12177 -26970
rect 12265 -27079 12286 -26970
rect 10553 -27084 12286 -27079
rect -30288 -30641 -27949 -30636
rect -30288 -30751 -30274 -30641
rect -30182 -30751 -27949 -30641
rect -30288 -30756 -27949 -30751
rect 10506 -30642 13923 -30636
rect 10506 -30751 13814 -30642
rect 13902 -30751 13923 -30642
rect 10506 -30756 13923 -30751
rect -30578 -34313 -27956 -34308
rect -30578 -34423 -30564 -34313
rect -30472 -34423 -27956 -34313
rect -30578 -34428 -27956 -34423
rect 10529 -34314 15558 -34308
rect 10529 -34423 15449 -34314
rect 15537 -34423 15558 -34314
rect 10529 -34428 15558 -34423
rect -30868 -37985 -27914 -37980
rect -30868 -38095 -30854 -37985
rect -30762 -38095 -27914 -37985
rect -30868 -38100 -27914 -38095
rect 10529 -37986 17195 -37980
rect 10529 -38095 17086 -37986
rect 17174 -38095 17195 -37986
rect 10529 -38100 17195 -38095
rect -31158 -41657 -27949 -41652
rect -31158 -41767 -31144 -41657
rect -31052 -41767 -27949 -41657
rect -31158 -41772 -27949 -41767
rect 10518 -41658 18830 -41652
rect 10518 -41767 18721 -41658
rect 18809 -41767 18830 -41658
rect 10518 -41772 18830 -41767
rect -31448 -45329 -27956 -45324
rect -31448 -45439 -31434 -45329
rect -31342 -45439 -27956 -45329
rect -31448 -45444 -27956 -45439
rect 10506 -45330 20466 -45324
rect 10506 -45439 20357 -45330
rect 20445 -45439 20466 -45330
rect 10506 -45444 20466 -45439
rect -31738 -49001 -27956 -48996
rect -31738 -49111 -31724 -49001
rect -31632 -49111 -27956 -49001
rect -31738 -49116 -27956 -49111
rect 10553 -49002 22103 -48996
rect 10553 -49111 21994 -49002
rect 22082 -49111 22103 -49002
rect 10553 -49116 22103 -49111
rect -32028 -52673 -27956 -52668
rect -32028 -52783 -32014 -52673
rect -31922 -52783 -27956 -52673
rect -32028 -52788 -27956 -52783
rect 10506 -52674 23739 -52668
rect 10506 -52783 23630 -52674
rect 23718 -52783 23739 -52674
rect 10506 -52788 23739 -52783
rect -4627 -54901 -4517 -54896
rect -4627 -55001 -4622 -54901
rect -4522 -55001 -4517 -54901
rect -4627 -55006 -4517 -55001
rect -1865 -54900 -1755 -54895
rect -1865 -55000 -1860 -54900
rect -1760 -55000 -1755 -54900
rect -1865 -55005 -1755 -55000
rect 894 -54899 1004 -54894
rect 894 -54999 899 -54899
rect 999 -54999 1004 -54899
rect 894 -55004 1004 -54999
rect 3654 -54900 3764 -54895
rect 3654 -55000 3659 -54900
rect 3759 -55000 3764 -54900
rect -4622 -58300 -4522 -55006
rect -1860 -58300 -1760 -55005
rect 899 -58300 999 -55004
rect 3654 -55005 3764 -55000
rect 6414 -54900 6524 -54895
rect 6414 -55000 6419 -54900
rect 6519 -55000 6524 -54900
rect 6414 -55005 6524 -55000
rect 9174 -54900 9284 -54895
rect 9174 -55000 9179 -54900
rect 9279 -55000 9284 -54900
rect 9174 -55005 9284 -55000
rect 3659 -58300 3759 -55005
rect 6419 -58300 6519 -55005
rect 9179 -58300 9279 -55005
<< via3 >>
rect 9338 13130 9648 13135
rect 9338 12835 9343 13130
rect 9343 12835 9643 13130
rect 9643 12835 9648 13130
rect 9342 11961 9642 12261
rect -12681 10599 -12381 10899
rect -11807 10899 -11507 10904
rect -11807 10599 -11512 10899
rect -11512 10599 -11507 10899
rect -11807 10594 -11507 10599
rect -2453 10528 -2153 10533
rect -2453 10228 -2158 10528
rect -2158 10228 -2153 10528
rect -2453 10223 -2153 10228
rect -2458 9687 -2158 9987
rect 850 10539 1451 10544
rect 850 9938 855 10539
rect 855 9938 1451 10539
rect 850 9933 1451 9938
rect 9056 10534 9657 10539
rect 9056 9933 9652 10534
rect 9652 9933 9657 10534
rect 9056 9928 9657 9933
rect 11563 10528 11863 10533
rect 11563 10228 11568 10528
rect 11568 10228 11863 10528
rect 11563 10223 11863 10228
rect 1633 9755 2234 9760
rect 1633 9154 2229 9755
rect 2229 9154 2234 9755
rect 1633 9149 2234 9154
rect 8300 9768 8901 9773
rect 8300 9167 8305 9768
rect 8305 9167 8901 9768
rect 11568 9687 11868 9987
rect 8300 9162 8901 9167
rect -21659 7791 -21359 8091
rect -20620 6296 -20320 6301
rect -20620 5996 -20615 6296
rect -20615 5996 -20320 6296
rect -20620 5991 -20320 5996
rect -45460 -6464 -45028 -6032
rect -15141 8701 -14841 8706
rect -19720 8331 -19715 8626
rect -19715 8331 -19415 8626
rect -19415 8331 -19410 8626
rect -15141 8401 -14846 8701
rect -14846 8401 -14841 8701
rect -15141 8396 -14841 8401
rect -19720 8326 -19410 8331
rect -13588 8122 -13288 8422
rect -15992 6659 -15692 6959
rect -18733 5460 -18433 5760
rect -11805 3340 -11495 3345
rect -15363 2903 -15063 3203
rect -11805 3045 -11800 3340
rect -11800 3045 -11500 3340
rect -11500 3045 -11495 3340
rect -16847 2298 -16537 2303
rect -16847 2003 -16842 2298
rect -16842 2003 -16542 2298
rect -16542 2003 -16537 2298
rect 8298 4336 8899 4341
rect 1637 4326 2238 4331
rect -2589 3794 -2584 4089
rect -2584 3794 -2284 4089
rect -2284 3794 -2279 4089
rect -2589 3789 -2279 3794
rect -1720 3794 -1715 4089
rect -1715 3794 -1415 4089
rect -1415 3794 -1410 4089
rect -1720 3789 -1410 3794
rect 1637 3725 2233 4326
rect 2233 3725 2238 4326
rect 1637 3720 2238 3725
rect 8298 3735 8894 4336
rect 8894 3735 8899 4336
rect 8298 3730 8899 3735
rect 883 3584 1484 3589
rect 883 2983 1479 3584
rect 1479 2983 1484 3584
rect 883 2978 1484 2983
rect 9080 3552 9681 3557
rect 9080 2951 9676 3552
rect 9676 2951 9681 3552
rect 9080 2946 9681 2951
rect -2855 2139 -2423 2144
rect -2855 1707 -2428 2139
rect -2428 1707 -2423 2139
rect -2855 1702 -2423 1707
rect 10869 2346 11169 2646
rect 11733 2346 11738 2641
rect 11738 2346 12038 2641
rect 12038 2346 12043 2641
rect 11733 2341 12043 2346
rect 5112 -932 5422 -927
rect 5112 -1227 5117 -932
rect 5117 -1227 5417 -932
rect 5417 -1227 5422 -932
rect 5117 -4687 5417 -4387
rect 25178 -6444 25610 -6012
rect 25531 -12795 25841 -12790
rect 25531 -13090 25536 -12795
rect 25536 -13090 25836 -12795
rect 25836 -13090 25841 -12795
rect 24527 -17054 24827 -16754
rect 26543 -17054 26843 -16754
<< metal4 >>
rect -54600 85800 39000 93800
rect -54600 14600 -46600 85800
rect -40153 66060 24652 72145
rect 23790 66044 24652 66060
rect -40176 27837 24573 33922
rect 23786 27818 24573 27837
rect 31000 14600 39000 85800
rect -54600 13135 39000 14600
rect -54600 12835 9338 13135
rect 9648 12835 39000 13135
rect -54600 12603 39000 12835
rect -54600 -2805 -52539 12603
rect -46169 -2805 -44415 12603
rect -54600 -2893 -44415 -2805
rect -22171 12544 39000 12603
rect -22171 12418 15667 12544
rect -22171 11808 9179 12418
rect 9303 12261 9671 12295
rect 9303 11961 9342 12261
rect 9642 11961 9671 12261
rect 9303 11927 9671 11961
rect 9789 11808 15667 12418
rect -22171 11250 15667 11808
rect -22171 11058 2807 11250
rect -22171 10448 -12836 11058
rect -12715 10899 -12347 10938
rect -12715 10599 -12681 10899
rect -12381 10599 -12347 10899
rect -12715 10570 -12347 10599
rect -12226 10904 2807 11058
rect -12226 10594 -11807 10904
rect -11507 10594 2807 10904
rect -12226 10544 2807 10594
rect -12226 10533 850 10544
rect -12226 10448 -2453 10533
rect -22171 10223 -2453 10448
rect -2153 10223 850 10533
rect -22171 10148 850 10223
rect -22171 9538 -2607 10148
rect -2487 9987 -2119 10021
rect -2487 9687 -2458 9987
rect -2158 9687 -2119 9987
rect -2487 9653 -2119 9687
rect -1997 9933 850 10148
rect 1451 9933 2807 10544
rect -1997 9893 2807 9933
rect 7724 10539 15667 11250
rect 7724 9928 9056 10539
rect 9657 10533 15667 10539
rect 9657 10223 11563 10533
rect 11863 10223 15667 10533
rect 9657 10151 15667 10223
rect 9657 9928 11409 10151
rect 7724 9893 11409 9928
rect -1997 9538 1534 9893
rect 8900 9773 8902 9774
rect -22171 8706 1534 9538
rect 1632 9760 1634 9761
rect 1632 9149 1633 9760
rect 8901 9162 8902 9773
rect 8900 9161 8902 9162
rect 8983 9541 11409 9893
rect 11529 9987 11897 10021
rect 11529 9687 11568 9987
rect 11868 9687 11897 9987
rect 11529 9653 11897 9687
rect 12019 9541 15667 10151
rect 1632 9148 1634 9149
rect -22171 8626 -15141 8706
rect -22171 8326 -19720 8626
rect -19410 8396 -15141 8626
rect -14841 8584 1534 8706
rect -14841 8396 -13744 8584
rect -19410 8326 -13744 8396
rect -22171 8269 -13744 8326
rect -22171 7659 -21813 8269
rect -21698 8091 -21330 8125
rect -21698 7791 -21659 8091
rect -21359 7791 -21330 8091
rect -21698 7757 -21330 7791
rect -21203 7974 -13744 8269
rect -13622 8422 -13254 8461
rect -13622 8122 -13588 8422
rect -13288 8122 -13254 8422
rect -13622 8093 -13254 8122
rect -13134 7974 1534 8584
rect -21203 7659 1534 7974
rect -22171 7120 1534 7659
rect -22171 6510 -16143 7120
rect -16021 6959 -15653 6993
rect -16021 6659 -15992 6959
rect -15692 6659 -15653 6959
rect -16021 6625 -15653 6659
rect -15533 6510 1534 7120
rect -22171 6301 1534 6510
rect -22171 5991 -20620 6301
rect -20320 5991 1534 6301
rect -22171 5943 1534 5991
rect -22171 5929 -18207 5943
rect -22171 5319 -18891 5929
rect -18767 5760 -18399 5789
rect -18767 5460 -18733 5760
rect -18433 5460 -18399 5760
rect -18767 5421 -18399 5460
rect -18281 5319 -18207 5929
rect -22171 3571 -18207 5319
rect -14389 4247 1534 5943
rect 8297 4341 8299 4342
rect -14389 3639 -2737 4247
rect -2125 4089 1534 4247
rect -2125 3789 -1720 4089
rect -1410 3789 1534 4089
rect -2125 3639 1534 3789
rect 1636 4331 1638 4332
rect 1636 3720 1637 4331
rect 8297 3730 8298 4341
rect 8297 3729 8299 3730
rect 1636 3719 1638 3720
rect 8983 3639 15667 9541
rect -14389 3589 2807 3639
rect -14389 3571 883 3589
rect -22171 3387 883 3571
rect -22171 2777 -15513 3387
rect -14903 3345 883 3387
rect -15402 3203 -15034 3237
rect -15402 2903 -15363 3203
rect -15063 2903 -15034 3203
rect -15402 2869 -15034 2903
rect -14903 3045 -11805 3345
rect -11495 3045 883 3345
rect -14903 2978 883 3045
rect 1484 2978 2807 3589
rect -14903 2777 2807 2978
rect -22171 2314 2807 2777
rect -22171 2303 -3008 2314
rect -22171 2003 -16847 2303
rect -16537 2003 -3008 2303
rect -2270 2292 2807 2314
rect 7724 3557 15667 3639
rect 7724 2946 9080 3557
rect 9681 2946 15667 3557
rect 7724 2802 15667 2946
rect 7724 2292 10706 2802
rect 10835 2646 11203 2675
rect 10835 2346 10869 2646
rect 11169 2346 11203 2646
rect 10835 2307 11203 2346
rect 11316 2641 15667 2802
rect 11316 2341 11733 2641
rect 12043 2341 15667 2641
rect -2270 2192 10706 2292
rect 11316 2192 15667 2341
rect -22171 1560 -3008 2003
rect -2856 2144 -2854 2145
rect -2856 1702 -2855 2144
rect -2856 1701 -2854 1702
rect -2270 1560 15667 2192
rect -22171 -927 15667 1560
rect -22171 -1227 5112 -927
rect 5422 -1227 15667 -927
rect -22171 -2890 15667 -1227
rect 23952 -2890 26008 12544
rect -22171 -2893 26008 -2890
rect -54600 -2914 26008 -2893
rect 36280 -2914 39000 12544
rect -54600 -4228 39000 -2914
rect -54600 -4838 4964 -4228
rect 5083 -4387 5451 -4358
rect 5083 -4687 5117 -4387
rect 5417 -4687 5451 -4387
rect 5083 -4726 5451 -4687
rect 5574 -4838 39000 -4228
rect -54600 -4881 39000 -4838
rect -54600 -4919 25967 -4881
rect -54600 -10212 -52480 -4919
rect -46260 -4927 25967 -4919
rect -46260 -5916 -44256 -4927
rect -46260 -6578 -45575 -5916
rect -45490 -6032 -45001 -6002
rect -45490 -6464 -45460 -6032
rect -45028 -6464 -45001 -6032
rect -45490 -6494 -45001 -6464
rect -44921 -6578 -44256 -5916
rect -46260 -10146 -44256 -6578
rect 24377 -5876 25967 -4927
rect 24377 -6567 25055 -5876
rect 25151 -6012 25640 -5982
rect 25151 -6444 25178 -6012
rect 25610 -6444 25640 -6012
rect 25151 -6474 25640 -6444
rect 25741 -6567 25967 -5876
rect 24377 -10146 25967 -6567
rect -46260 -10210 25967 -10146
rect 36507 -10210 39000 -4881
rect -46260 -10212 39000 -10210
rect -54600 -12790 39000 -10212
rect -54600 -13090 25531 -12790
rect 25841 -13090 39000 -12790
rect -54600 -13782 39000 -13090
rect -54600 -54681 -52378 -13782
rect -30786 -13788 39000 -13782
rect -30786 -13800 27250 -13788
rect -30786 -54681 -28200 -13800
rect -23868 -16428 -23548 -13800
rect 6852 -16428 7172 -13800
rect 10600 -13823 27250 -13800
rect 10600 -17604 12914 -13823
rect 24135 -16592 27250 -13823
rect 24135 -17202 24384 -16592
rect 24994 -16593 27250 -16592
rect 24498 -16753 24866 -16720
rect 24498 -17057 24527 -16753
rect 24831 -17057 24866 -16753
rect 24498 -17088 24866 -17057
rect 24994 -17202 26373 -16593
rect 26504 -16752 26872 -16720
rect 26504 -17055 26541 -16752
rect 26847 -17055 26872 -16752
rect 26504 -17088 26872 -17055
rect 24135 -17203 26373 -17202
rect 26983 -17203 27250 -16593
rect 24135 -17588 27250 -17203
rect 36510 -17604 39000 -13788
rect -54600 -54800 -28200 -54681
rect -23868 -54800 -23548 -52202
rect 6852 -54800 7172 -52116
rect 10600 -54681 12951 -17604
rect 36411 -54681 39000 -17604
rect 10600 -54800 39000 -54681
rect -54600 -58200 39000 -54800
<< via4 >>
rect -46238 66060 -40153 72145
rect 24652 66044 30624 72129
rect -46261 27837 -40176 33922
rect 24573 27818 30620 33903
rect 9342 11961 9642 12261
rect -12681 10599 -12381 10899
rect -2458 9687 -2158 9987
rect 8299 9773 8900 9774
rect 1634 9760 2235 9761
rect 1634 9149 2234 9760
rect 2234 9149 2235 9760
rect 8299 9162 8300 9773
rect 8300 9162 8900 9773
rect 8299 9161 8900 9162
rect 11568 9687 11868 9987
rect 1634 9148 2235 9149
rect -21659 7791 -21359 8091
rect -13588 8122 -13288 8422
rect -15992 6659 -15692 6959
rect -18733 5460 -18433 5760
rect 8299 4341 8900 4342
rect -2594 4089 -2274 4099
rect -2594 3789 -2589 4089
rect -2589 3789 -2279 4089
rect -2279 3789 -2274 4089
rect -2594 3779 -2274 3789
rect 1638 4331 2239 4332
rect 1638 3720 2238 4331
rect 2238 3720 2239 4331
rect 8299 3730 8899 4341
rect 8899 3730 8900 4341
rect 8299 3729 8900 3730
rect 1638 3719 2239 3720
rect -15363 2903 -15063 3203
rect 10869 2346 11169 2646
rect -2854 2144 -2422 2145
rect -2854 1702 -2423 2144
rect -2423 1702 -2422 2144
rect -2854 1701 -2422 1702
rect 5117 -4687 5417 -4387
rect -45460 -6464 -45028 -6032
rect 25178 -6444 25610 -6012
rect 24527 -16754 24831 -16753
rect 24527 -17054 24827 -16754
rect 24827 -17054 24831 -16754
rect 24527 -17057 24831 -17054
rect 26541 -16754 26847 -16752
rect 26541 -17054 26543 -16754
rect 26543 -17054 26843 -16754
rect 26843 -17054 26847 -16754
rect 26541 -17055 26847 -17054
<< metal5 >>
rect -54600 83954 39000 93800
rect -54600 72145 -38820 83954
rect -54600 66060 -46238 72145
rect -40153 66060 -38820 72145
rect -54600 33922 -38820 66060
rect -54600 27837 -46261 33922
rect -40176 27837 -38820 33922
rect -54600 15907 -38820 27837
rect 22834 72129 39000 83954
rect 22834 66044 24652 72129
rect 30624 66044 39000 72129
rect 22834 33903 39000 66044
rect 22834 27818 24573 33903
rect 30620 27818 39000 33903
rect 22834 15907 39000 27818
rect -54600 14732 39000 15907
rect -54600 -2814 -52496 14732
rect -46236 13381 26034 14732
rect -46236 13226 15686 13381
rect -46236 -2814 -44330 13226
rect -54600 -2945 -44330 -2814
rect -22252 12261 15686 13226
rect -22252 11961 9342 12261
rect 9642 11961 15686 12261
rect -22252 10899 15686 11961
rect -22252 10599 -12681 10899
rect -12381 10599 15686 10899
rect -22252 9987 15686 10599
rect -22252 9687 -2458 9987
rect -2158 9774 11568 9987
rect -2158 9761 8299 9774
rect -2158 9687 1634 9761
rect -22252 9148 1634 9687
rect 2235 9161 8299 9761
rect 8900 9687 11568 9774
rect 11868 9687 15686 9987
rect 8900 9161 15686 9687
rect 2235 9148 15686 9161
rect -22252 8422 15686 9148
rect -22252 8122 -13588 8422
rect -13288 8122 15686 8422
rect -22252 8091 15686 8122
rect -22252 7791 -21659 8091
rect -21359 7791 15686 8091
rect -22252 6959 15686 7791
rect -22252 6659 -15992 6959
rect -15692 6659 15686 6959
rect -22252 5760 15686 6659
rect -22252 5460 -18733 5760
rect -18433 5460 15686 5760
rect -22252 4342 15686 5460
rect -22252 4332 8299 4342
rect -22252 4099 1638 4332
rect -22252 3779 -2594 4099
rect -2274 3779 1638 4099
rect -22252 3719 1638 3779
rect 2239 3729 8299 4332
rect 8900 3729 15686 4342
rect 2239 3719 15686 3729
rect -22252 3203 15686 3719
rect -22252 2903 -15363 3203
rect -15063 2903 15686 3203
rect -22252 2646 15686 2903
rect -22252 2346 10869 2646
rect 11169 2346 15686 2646
rect -22252 2145 15686 2346
rect -22252 1701 -2854 2145
rect -2422 1701 15686 2145
rect -22252 -2867 15686 1701
rect 23927 -2867 26034 13381
rect -22252 -2908 26034 -2867
rect 36277 -2908 39000 14732
rect -22252 -2945 39000 -2908
rect -54600 -4387 39000 -2945
rect -54600 -4687 5117 -4387
rect 5417 -4687 39000 -4387
rect -54600 -4879 39000 -4687
rect -54600 -4928 26027 -4879
rect -54600 -10194 -52480 -4928
rect -46287 -6032 -44239 -4928
rect -46287 -6464 -45460 -6032
rect -45028 -6464 -44239 -6032
rect -46287 -10146 -44239 -6464
rect 24369 -6012 26027 -4928
rect 24369 -6444 25178 -6012
rect 25610 -6444 26027 -6012
rect 24369 -10146 26027 -6444
rect -46287 -10194 26027 -10146
rect 36462 -10194 39000 -4879
rect -54600 -13841 39000 -10194
rect -54600 -13864 12972 -13841
rect -54600 -13938 -28076 -13864
rect -54600 -54619 -52370 -13938
rect -30816 -17738 -28076 -13938
rect 10562 -17738 12972 -13864
rect 24093 -16752 27290 -13841
rect 24093 -16753 26541 -16752
rect 24093 -17057 24527 -16753
rect 24831 -17055 26541 -16753
rect 26847 -17055 27290 -16752
rect 24831 -17057 27290 -17055
rect 24093 -17530 27290 -17057
rect -30816 -18058 -26700 -17738
rect 9280 -18058 12972 -17738
rect -30816 -48374 -28076 -18058
rect 10562 -48374 12972 -18058
rect -30816 -48694 -26700 -48374
rect 9280 -48694 12972 -48374
rect -30816 -54619 -28076 -48694
rect -54600 -54700 -28076 -54619
rect 10562 -54619 12972 -48694
rect 36468 -54619 39000 -13841
rect 10562 -54700 39000 -54619
rect -54600 -58300 39000 -54700
use full_vco_1  full_vco_1_0
timestamp 1669280253
transform 1 0 1247 0 1 3352
box -7141 -8039 14057 8505
use inv_buffer2  inv_buffer2_0
timestamp 1668357910
transform 0 1 24547 1 0 -16070
box 0 0 2204 1138
use inv_buffer2  inv_buffer2_1
timestamp 1668357910
transform 0 -1 26823 1 0 -16070
box 0 0 2204 1138
use inv_buffer2  inv_buffer2_8
timestamp 1668357910
transform 0 1 -21233 -1 0 8898
box 0 0 2204 1138
use inv_buffer2  inv_buffer2_9
timestamp 1668357910
transform -1 0 12197 0 1 11981
box 0 0 2204 1138
use r2r_8  r2r_8_0
timestamp 1668357910
transform -1 0 25125 0 1 -10561
box -485 -593 13937 10023
use r2r_8  r2r_8_1
timestamp 1668357910
transform 1 0 -30985 0 1 -10581
box -485 -593 13937 10023
use r2r_8  r2r_8_2
timestamp 1668357910
transform 1 0 -44975 0 1 -10581
box -485 -593 13937 10023
use r2r_10  r2r_10_0
timestamp 1668357910
transform 1 0 -16995 0 1 -10581
box -485 -593 17209 10023
use slopebuf  slopebuf_0
timestamp 1669280253
transform 1 0 -19311 0 1 6012
box -866 -1740 4686 2950
use sspd  sspd_0
timestamp 1669280253
transform 0 1 -16419 -1 0 9251
box -1125 214 7472 5865
use voltage_control  voltage_control_0
timestamp 1669279853
transform 1 0 -80552 0 1 -4512
box 41052 6053 104762 89673
<< labels >>
rlabel via2 9343 12830 9643 13130 0 vdd
port 1 n
rlabel via2 -45460 -6464 -45028 -6032 6 vss
rlabel via2 25178 -6444 25610 -6012 5 vss
rlabel via2 24527 -17054 24827 -16754 0 vss
rlabel via2 26543 -17054 26843 -16754 3 vss
rlabel via2 25536 -13095 25836 -12795 2 vdd
rlabel via2 10869 2346 11169 2646 0 vss
rlabel via2 11738 2346 12038 2646 0 vdd
rlabel via2 -11812 10599 -11512 10899 4 vdd
rlabel via2 -11800 3040 -11500 3340 0 vdd
rlabel via2 -16842 1998 -16542 2298 0 vdd
rlabel via2 -12681 10599 -12381 10899 5 vss
rlabel via2 -13588 8122 -13288 8422 0 vss
rlabel via2 -15146 8401 -14846 8701 6 vdd
rlabel via2 -18733 5460 -18433 5760 7 vss
rlabel via2 -19715 8331 -19415 8631 0 vdd
rlabel via2 -15992 6659 -15692 6959 3 vss
rlabel via2 -21659 7791 -21359 8091 0 vss
rlabel via2 -20615 5996 -20315 6296 0 vdd
rlabel via1 855 9938 1456 10539 0 vdd
rlabel metal1 8304 9167 8905 9768 7 vss
rlabel metal4 -11042 27837 -4877 33922 7 vss
rlabel metal4 -11042 66060 -4877 72145 7 vss
rlabel via2 9342 11961 9642 12261 0 vss
port 2 n
rlabel metal1 1626 3725 2227 4326 0 vss
rlabel metal1 1622 9154 2223 9755 0 vss
rlabel metal1 8287 3735 8888 4336 0 vss
rlabel via1 9075 2951 9676 3552 5 vdd
rlabel via1 9051 9933 9652 10534 5 vdd
rlabel via1 878 2983 1479 3584 5 vdd
rlabel via2 -15363 2903 -15063 3203 0 vss
rlabel metal3 -4622 -58298 -4522 -58198 6 reset
port 3 n
rlabel metal3 -1860 -58300 -1760 -58200 3 clk_in
port 4 n
rlabel metal3 899 -58300 999 -58200 7 read
port 5 n
rlabel metal3 3659 -58282 3759 -58182 0 load
port 6 n
rlabel metal3 6419 -58282 6519 -58182 5 s_in
port 7 n
rlabel metal3 9179 -58282 9279 -58182 0 s_out
port 8 n
rlabel metal1 25632 -16189 25752 -16069 6 ref_in
port 9 n
rlabel metal1 14915 9152 14955 9192 8 out
port 10 n
rlabel metal2 25008 -13720 25128 -13600 0 ref_digital
rlabel metal3 -1081 -403 -1015 -337 0 vcoarse
rlabel metal3 682 -421 748 -355 7 lock
<< end >>
