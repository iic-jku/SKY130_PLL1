magic
tech sky130A
magscale 1 2
timestamp 1662021593
<< viali >>
rect 1409 7361 1443 7395
rect 5825 4981 5859 5015
<< metal1 >>
rect 1104 7642 6532 7664
rect 1104 7590 2759 7642
rect 2811 7590 2823 7642
rect 2875 7590 2887 7642
rect 2939 7590 2951 7642
rect 3003 7590 3015 7642
rect 3067 7590 4568 7642
rect 4620 7590 4632 7642
rect 4684 7590 4696 7642
rect 4748 7590 4760 7642
rect 4812 7590 4824 7642
rect 4876 7590 6532 7642
rect 1104 7568 6532 7590
rect 1394 7392 1400 7404
rect 1355 7364 1400 7392
rect 1394 7352 1400 7364
rect 1452 7352 1458 7404
rect 1104 7098 6532 7120
rect 1104 7046 1854 7098
rect 1906 7046 1918 7098
rect 1970 7046 1982 7098
rect 2034 7046 2046 7098
rect 2098 7046 2110 7098
rect 2162 7046 3664 7098
rect 3716 7046 3728 7098
rect 3780 7046 3792 7098
rect 3844 7046 3856 7098
rect 3908 7046 3920 7098
rect 3972 7046 5473 7098
rect 5525 7046 5537 7098
rect 5589 7046 5601 7098
rect 5653 7046 5665 7098
rect 5717 7046 5729 7098
rect 5781 7046 6532 7098
rect 1104 7024 6532 7046
rect 1104 6554 6532 6576
rect 1104 6502 2759 6554
rect 2811 6502 2823 6554
rect 2875 6502 2887 6554
rect 2939 6502 2951 6554
rect 3003 6502 3015 6554
rect 3067 6502 4568 6554
rect 4620 6502 4632 6554
rect 4684 6502 4696 6554
rect 4748 6502 4760 6554
rect 4812 6502 4824 6554
rect 4876 6502 6532 6554
rect 1104 6480 6532 6502
rect 1104 6010 6532 6032
rect 1104 5958 1854 6010
rect 1906 5958 1918 6010
rect 1970 5958 1982 6010
rect 2034 5958 2046 6010
rect 2098 5958 2110 6010
rect 2162 5958 3664 6010
rect 3716 5958 3728 6010
rect 3780 5958 3792 6010
rect 3844 5958 3856 6010
rect 3908 5958 3920 6010
rect 3972 5958 5473 6010
rect 5525 5958 5537 6010
rect 5589 5958 5601 6010
rect 5653 5958 5665 6010
rect 5717 5958 5729 6010
rect 5781 5958 6532 6010
rect 1104 5936 6532 5958
rect 1104 5466 6532 5488
rect 1104 5414 2759 5466
rect 2811 5414 2823 5466
rect 2875 5414 2887 5466
rect 2939 5414 2951 5466
rect 3003 5414 3015 5466
rect 3067 5414 4568 5466
rect 4620 5414 4632 5466
rect 4684 5414 4696 5466
rect 4748 5414 4760 5466
rect 4812 5414 4824 5466
rect 4876 5414 6532 5466
rect 1104 5392 6532 5414
rect 5813 5015 5871 5021
rect 5813 4981 5825 5015
rect 5859 5012 5871 5015
rect 5902 5012 5908 5024
rect 5859 4984 5908 5012
rect 5859 4981 5871 4984
rect 5813 4975 5871 4981
rect 5902 4972 5908 4984
rect 5960 4972 5966 5024
rect 1104 4922 6532 4944
rect 1104 4870 1854 4922
rect 1906 4870 1918 4922
rect 1970 4870 1982 4922
rect 2034 4870 2046 4922
rect 2098 4870 2110 4922
rect 2162 4870 3664 4922
rect 3716 4870 3728 4922
rect 3780 4870 3792 4922
rect 3844 4870 3856 4922
rect 3908 4870 3920 4922
rect 3972 4870 5473 4922
rect 5525 4870 5537 4922
rect 5589 4870 5601 4922
rect 5653 4870 5665 4922
rect 5717 4870 5729 4922
rect 5781 4870 6532 4922
rect 1104 4848 6532 4870
rect 1104 4378 6532 4400
rect 1104 4326 2759 4378
rect 2811 4326 2823 4378
rect 2875 4326 2887 4378
rect 2939 4326 2951 4378
rect 3003 4326 3015 4378
rect 3067 4326 4568 4378
rect 4620 4326 4632 4378
rect 4684 4326 4696 4378
rect 4748 4326 4760 4378
rect 4812 4326 4824 4378
rect 4876 4326 6532 4378
rect 1104 4304 6532 4326
rect 1104 3834 6532 3856
rect 1104 3782 1854 3834
rect 1906 3782 1918 3834
rect 1970 3782 1982 3834
rect 2034 3782 2046 3834
rect 2098 3782 2110 3834
rect 2162 3782 3664 3834
rect 3716 3782 3728 3834
rect 3780 3782 3792 3834
rect 3844 3782 3856 3834
rect 3908 3782 3920 3834
rect 3972 3782 5473 3834
rect 5525 3782 5537 3834
rect 5589 3782 5601 3834
rect 5653 3782 5665 3834
rect 5717 3782 5729 3834
rect 5781 3782 6532 3834
rect 1104 3760 6532 3782
rect 1104 3290 6532 3312
rect 1104 3238 2759 3290
rect 2811 3238 2823 3290
rect 2875 3238 2887 3290
rect 2939 3238 2951 3290
rect 3003 3238 3015 3290
rect 3067 3238 4568 3290
rect 4620 3238 4632 3290
rect 4684 3238 4696 3290
rect 4748 3238 4760 3290
rect 4812 3238 4824 3290
rect 4876 3238 6532 3290
rect 1104 3216 6532 3238
rect 1104 2746 6532 2768
rect 1104 2694 1854 2746
rect 1906 2694 1918 2746
rect 1970 2694 1982 2746
rect 2034 2694 2046 2746
rect 2098 2694 2110 2746
rect 2162 2694 3664 2746
rect 3716 2694 3728 2746
rect 3780 2694 3792 2746
rect 3844 2694 3856 2746
rect 3908 2694 3920 2746
rect 3972 2694 5473 2746
rect 5525 2694 5537 2746
rect 5589 2694 5601 2746
rect 5653 2694 5665 2746
rect 5717 2694 5729 2746
rect 5781 2694 6532 2746
rect 1104 2672 6532 2694
rect 1104 2202 6532 2224
rect 1104 2150 2759 2202
rect 2811 2150 2823 2202
rect 2875 2150 2887 2202
rect 2939 2150 2951 2202
rect 3003 2150 3015 2202
rect 3067 2150 4568 2202
rect 4620 2150 4632 2202
rect 4684 2150 4696 2202
rect 4748 2150 4760 2202
rect 4812 2150 4824 2202
rect 4876 2150 6532 2202
rect 1104 2128 6532 2150
<< via1 >>
rect 2759 7590 2811 7642
rect 2823 7590 2875 7642
rect 2887 7590 2939 7642
rect 2951 7590 3003 7642
rect 3015 7590 3067 7642
rect 4568 7590 4620 7642
rect 4632 7590 4684 7642
rect 4696 7590 4748 7642
rect 4760 7590 4812 7642
rect 4824 7590 4876 7642
rect 1400 7395 1452 7404
rect 1400 7361 1409 7395
rect 1409 7361 1443 7395
rect 1443 7361 1452 7395
rect 1400 7352 1452 7361
rect 1854 7046 1906 7098
rect 1918 7046 1970 7098
rect 1982 7046 2034 7098
rect 2046 7046 2098 7098
rect 2110 7046 2162 7098
rect 3664 7046 3716 7098
rect 3728 7046 3780 7098
rect 3792 7046 3844 7098
rect 3856 7046 3908 7098
rect 3920 7046 3972 7098
rect 5473 7046 5525 7098
rect 5537 7046 5589 7098
rect 5601 7046 5653 7098
rect 5665 7046 5717 7098
rect 5729 7046 5781 7098
rect 2759 6502 2811 6554
rect 2823 6502 2875 6554
rect 2887 6502 2939 6554
rect 2951 6502 3003 6554
rect 3015 6502 3067 6554
rect 4568 6502 4620 6554
rect 4632 6502 4684 6554
rect 4696 6502 4748 6554
rect 4760 6502 4812 6554
rect 4824 6502 4876 6554
rect 1854 5958 1906 6010
rect 1918 5958 1970 6010
rect 1982 5958 2034 6010
rect 2046 5958 2098 6010
rect 2110 5958 2162 6010
rect 3664 5958 3716 6010
rect 3728 5958 3780 6010
rect 3792 5958 3844 6010
rect 3856 5958 3908 6010
rect 3920 5958 3972 6010
rect 5473 5958 5525 6010
rect 5537 5958 5589 6010
rect 5601 5958 5653 6010
rect 5665 5958 5717 6010
rect 5729 5958 5781 6010
rect 2759 5414 2811 5466
rect 2823 5414 2875 5466
rect 2887 5414 2939 5466
rect 2951 5414 3003 5466
rect 3015 5414 3067 5466
rect 4568 5414 4620 5466
rect 4632 5414 4684 5466
rect 4696 5414 4748 5466
rect 4760 5414 4812 5466
rect 4824 5414 4876 5466
rect 5908 4972 5960 5024
rect 1854 4870 1906 4922
rect 1918 4870 1970 4922
rect 1982 4870 2034 4922
rect 2046 4870 2098 4922
rect 2110 4870 2162 4922
rect 3664 4870 3716 4922
rect 3728 4870 3780 4922
rect 3792 4870 3844 4922
rect 3856 4870 3908 4922
rect 3920 4870 3972 4922
rect 5473 4870 5525 4922
rect 5537 4870 5589 4922
rect 5601 4870 5653 4922
rect 5665 4870 5717 4922
rect 5729 4870 5781 4922
rect 2759 4326 2811 4378
rect 2823 4326 2875 4378
rect 2887 4326 2939 4378
rect 2951 4326 3003 4378
rect 3015 4326 3067 4378
rect 4568 4326 4620 4378
rect 4632 4326 4684 4378
rect 4696 4326 4748 4378
rect 4760 4326 4812 4378
rect 4824 4326 4876 4378
rect 1854 3782 1906 3834
rect 1918 3782 1970 3834
rect 1982 3782 2034 3834
rect 2046 3782 2098 3834
rect 2110 3782 2162 3834
rect 3664 3782 3716 3834
rect 3728 3782 3780 3834
rect 3792 3782 3844 3834
rect 3856 3782 3908 3834
rect 3920 3782 3972 3834
rect 5473 3782 5525 3834
rect 5537 3782 5589 3834
rect 5601 3782 5653 3834
rect 5665 3782 5717 3834
rect 5729 3782 5781 3834
rect 2759 3238 2811 3290
rect 2823 3238 2875 3290
rect 2887 3238 2939 3290
rect 2951 3238 3003 3290
rect 3015 3238 3067 3290
rect 4568 3238 4620 3290
rect 4632 3238 4684 3290
rect 4696 3238 4748 3290
rect 4760 3238 4812 3290
rect 4824 3238 4876 3290
rect 1854 2694 1906 2746
rect 1918 2694 1970 2746
rect 1982 2694 2034 2746
rect 2046 2694 2098 2746
rect 2110 2694 2162 2746
rect 3664 2694 3716 2746
rect 3728 2694 3780 2746
rect 3792 2694 3844 2746
rect 3856 2694 3908 2746
rect 3920 2694 3972 2746
rect 5473 2694 5525 2746
rect 5537 2694 5589 2746
rect 5601 2694 5653 2746
rect 5665 2694 5717 2746
rect 5729 2694 5781 2746
rect 2759 2150 2811 2202
rect 2823 2150 2875 2202
rect 2887 2150 2939 2202
rect 2951 2150 3003 2202
rect 3015 2150 3067 2202
rect 4568 2150 4620 2202
rect 4632 2150 4684 2202
rect 4696 2150 4748 2202
rect 4760 2150 4812 2202
rect 4824 2150 4876 2202
<< metal2 >>
rect 938 9194 994 9832
rect 938 9166 1348 9194
rect 938 9032 994 9166
rect 1320 8242 1348 9166
rect 2870 9032 2926 9832
rect 4802 9032 4858 9832
rect 6734 9032 6790 9832
rect 1320 8214 1440 8242
rect 1412 7410 1440 8214
rect 2759 7644 3067 7664
rect 2759 7642 2765 7644
rect 2821 7642 2845 7644
rect 2901 7642 2925 7644
rect 2981 7642 3005 7644
rect 3061 7642 3067 7644
rect 2821 7590 2823 7642
rect 3003 7590 3005 7642
rect 2759 7588 2765 7590
rect 2821 7588 2845 7590
rect 2901 7588 2925 7590
rect 2981 7588 3005 7590
rect 3061 7588 3067 7590
rect 2759 7568 3067 7588
rect 4568 7644 4876 7664
rect 4568 7642 4574 7644
rect 4630 7642 4654 7644
rect 4710 7642 4734 7644
rect 4790 7642 4814 7644
rect 4870 7642 4876 7644
rect 4630 7590 4632 7642
rect 4812 7590 4814 7642
rect 4568 7588 4574 7590
rect 4630 7588 4654 7590
rect 4710 7588 4734 7590
rect 4790 7588 4814 7590
rect 4870 7588 4876 7590
rect 4568 7568 4876 7588
rect 1400 7404 1452 7410
rect 1400 7346 1452 7352
rect 1854 7100 2162 7120
rect 1854 7098 1860 7100
rect 1916 7098 1940 7100
rect 1996 7098 2020 7100
rect 2076 7098 2100 7100
rect 2156 7098 2162 7100
rect 1916 7046 1918 7098
rect 2098 7046 2100 7098
rect 1854 7044 1860 7046
rect 1916 7044 1940 7046
rect 1996 7044 2020 7046
rect 2076 7044 2100 7046
rect 2156 7044 2162 7046
rect 1854 7024 2162 7044
rect 3664 7100 3972 7120
rect 3664 7098 3670 7100
rect 3726 7098 3750 7100
rect 3806 7098 3830 7100
rect 3886 7098 3910 7100
rect 3966 7098 3972 7100
rect 3726 7046 3728 7098
rect 3908 7046 3910 7098
rect 3664 7044 3670 7046
rect 3726 7044 3750 7046
rect 3806 7044 3830 7046
rect 3886 7044 3910 7046
rect 3966 7044 3972 7046
rect 3664 7024 3972 7044
rect 5473 7100 5781 7120
rect 5473 7098 5479 7100
rect 5535 7098 5559 7100
rect 5615 7098 5639 7100
rect 5695 7098 5719 7100
rect 5775 7098 5781 7100
rect 5535 7046 5537 7098
rect 5717 7046 5719 7098
rect 5473 7044 5479 7046
rect 5535 7044 5559 7046
rect 5615 7044 5639 7046
rect 5695 7044 5719 7046
rect 5775 7044 5781 7046
rect 5473 7024 5781 7044
rect 2759 6556 3067 6576
rect 2759 6554 2765 6556
rect 2821 6554 2845 6556
rect 2901 6554 2925 6556
rect 2981 6554 3005 6556
rect 3061 6554 3067 6556
rect 2821 6502 2823 6554
rect 3003 6502 3005 6554
rect 2759 6500 2765 6502
rect 2821 6500 2845 6502
rect 2901 6500 2925 6502
rect 2981 6500 3005 6502
rect 3061 6500 3067 6502
rect 2759 6480 3067 6500
rect 4568 6556 4876 6576
rect 4568 6554 4574 6556
rect 4630 6554 4654 6556
rect 4710 6554 4734 6556
rect 4790 6554 4814 6556
rect 4870 6554 4876 6556
rect 4630 6502 4632 6554
rect 4812 6502 4814 6554
rect 4568 6500 4574 6502
rect 4630 6500 4654 6502
rect 4710 6500 4734 6502
rect 4790 6500 4814 6502
rect 4870 6500 4876 6502
rect 4568 6480 4876 6500
rect 1854 6012 2162 6032
rect 1854 6010 1860 6012
rect 1916 6010 1940 6012
rect 1996 6010 2020 6012
rect 2076 6010 2100 6012
rect 2156 6010 2162 6012
rect 1916 5958 1918 6010
rect 2098 5958 2100 6010
rect 1854 5956 1860 5958
rect 1916 5956 1940 5958
rect 1996 5956 2020 5958
rect 2076 5956 2100 5958
rect 2156 5956 2162 5958
rect 1854 5936 2162 5956
rect 3664 6012 3972 6032
rect 3664 6010 3670 6012
rect 3726 6010 3750 6012
rect 3806 6010 3830 6012
rect 3886 6010 3910 6012
rect 3966 6010 3972 6012
rect 3726 5958 3728 6010
rect 3908 5958 3910 6010
rect 3664 5956 3670 5958
rect 3726 5956 3750 5958
rect 3806 5956 3830 5958
rect 3886 5956 3910 5958
rect 3966 5956 3972 5958
rect 3664 5936 3972 5956
rect 5473 6012 5781 6032
rect 5473 6010 5479 6012
rect 5535 6010 5559 6012
rect 5615 6010 5639 6012
rect 5695 6010 5719 6012
rect 5775 6010 5781 6012
rect 5535 5958 5537 6010
rect 5717 5958 5719 6010
rect 5473 5956 5479 5958
rect 5535 5956 5559 5958
rect 5615 5956 5639 5958
rect 5695 5956 5719 5958
rect 5775 5956 5781 5958
rect 5473 5936 5781 5956
rect 2759 5468 3067 5488
rect 2759 5466 2765 5468
rect 2821 5466 2845 5468
rect 2901 5466 2925 5468
rect 2981 5466 3005 5468
rect 3061 5466 3067 5468
rect 2821 5414 2823 5466
rect 3003 5414 3005 5466
rect 2759 5412 2765 5414
rect 2821 5412 2845 5414
rect 2901 5412 2925 5414
rect 2981 5412 3005 5414
rect 3061 5412 3067 5414
rect 2759 5392 3067 5412
rect 4568 5468 4876 5488
rect 4568 5466 4574 5468
rect 4630 5466 4654 5468
rect 4710 5466 4734 5468
rect 4790 5466 4814 5468
rect 4870 5466 4876 5468
rect 4630 5414 4632 5466
rect 4812 5414 4814 5466
rect 4568 5412 4574 5414
rect 4630 5412 4654 5414
rect 4710 5412 4734 5414
rect 4790 5412 4814 5414
rect 4870 5412 4876 5414
rect 4568 5392 4876 5412
rect 5908 5024 5960 5030
rect 5906 4992 5908 5001
rect 5960 4992 5962 5001
rect 1854 4924 2162 4944
rect 1854 4922 1860 4924
rect 1916 4922 1940 4924
rect 1996 4922 2020 4924
rect 2076 4922 2100 4924
rect 2156 4922 2162 4924
rect 1916 4870 1918 4922
rect 2098 4870 2100 4922
rect 1854 4868 1860 4870
rect 1916 4868 1940 4870
rect 1996 4868 2020 4870
rect 2076 4868 2100 4870
rect 2156 4868 2162 4870
rect 1854 4848 2162 4868
rect 3664 4924 3972 4944
rect 3664 4922 3670 4924
rect 3726 4922 3750 4924
rect 3806 4922 3830 4924
rect 3886 4922 3910 4924
rect 3966 4922 3972 4924
rect 3726 4870 3728 4922
rect 3908 4870 3910 4922
rect 3664 4868 3670 4870
rect 3726 4868 3750 4870
rect 3806 4868 3830 4870
rect 3886 4868 3910 4870
rect 3966 4868 3972 4870
rect 3664 4848 3972 4868
rect 5473 4924 5781 4944
rect 5906 4927 5962 4936
rect 5473 4922 5479 4924
rect 5535 4922 5559 4924
rect 5615 4922 5639 4924
rect 5695 4922 5719 4924
rect 5775 4922 5781 4924
rect 5535 4870 5537 4922
rect 5717 4870 5719 4922
rect 5473 4868 5479 4870
rect 5535 4868 5559 4870
rect 5615 4868 5639 4870
rect 5695 4868 5719 4870
rect 5775 4868 5781 4870
rect 5473 4848 5781 4868
rect 2759 4380 3067 4400
rect 2759 4378 2765 4380
rect 2821 4378 2845 4380
rect 2901 4378 2925 4380
rect 2981 4378 3005 4380
rect 3061 4378 3067 4380
rect 2821 4326 2823 4378
rect 3003 4326 3005 4378
rect 2759 4324 2765 4326
rect 2821 4324 2845 4326
rect 2901 4324 2925 4326
rect 2981 4324 3005 4326
rect 3061 4324 3067 4326
rect 2759 4304 3067 4324
rect 4568 4380 4876 4400
rect 4568 4378 4574 4380
rect 4630 4378 4654 4380
rect 4710 4378 4734 4380
rect 4790 4378 4814 4380
rect 4870 4378 4876 4380
rect 4630 4326 4632 4378
rect 4812 4326 4814 4378
rect 4568 4324 4574 4326
rect 4630 4324 4654 4326
rect 4710 4324 4734 4326
rect 4790 4324 4814 4326
rect 4870 4324 4876 4326
rect 4568 4304 4876 4324
rect 1854 3836 2162 3856
rect 1854 3834 1860 3836
rect 1916 3834 1940 3836
rect 1996 3834 2020 3836
rect 2076 3834 2100 3836
rect 2156 3834 2162 3836
rect 1916 3782 1918 3834
rect 2098 3782 2100 3834
rect 1854 3780 1860 3782
rect 1916 3780 1940 3782
rect 1996 3780 2020 3782
rect 2076 3780 2100 3782
rect 2156 3780 2162 3782
rect 1854 3760 2162 3780
rect 3664 3836 3972 3856
rect 3664 3834 3670 3836
rect 3726 3834 3750 3836
rect 3806 3834 3830 3836
rect 3886 3834 3910 3836
rect 3966 3834 3972 3836
rect 3726 3782 3728 3834
rect 3908 3782 3910 3834
rect 3664 3780 3670 3782
rect 3726 3780 3750 3782
rect 3806 3780 3830 3782
rect 3886 3780 3910 3782
rect 3966 3780 3972 3782
rect 3664 3760 3972 3780
rect 5473 3836 5781 3856
rect 5473 3834 5479 3836
rect 5535 3834 5559 3836
rect 5615 3834 5639 3836
rect 5695 3834 5719 3836
rect 5775 3834 5781 3836
rect 5535 3782 5537 3834
rect 5717 3782 5719 3834
rect 5473 3780 5479 3782
rect 5535 3780 5559 3782
rect 5615 3780 5639 3782
rect 5695 3780 5719 3782
rect 5775 3780 5781 3782
rect 5473 3760 5781 3780
rect 2759 3292 3067 3312
rect 2759 3290 2765 3292
rect 2821 3290 2845 3292
rect 2901 3290 2925 3292
rect 2981 3290 3005 3292
rect 3061 3290 3067 3292
rect 2821 3238 2823 3290
rect 3003 3238 3005 3290
rect 2759 3236 2765 3238
rect 2821 3236 2845 3238
rect 2901 3236 2925 3238
rect 2981 3236 3005 3238
rect 3061 3236 3067 3238
rect 2759 3216 3067 3236
rect 4568 3292 4876 3312
rect 4568 3290 4574 3292
rect 4630 3290 4654 3292
rect 4710 3290 4734 3292
rect 4790 3290 4814 3292
rect 4870 3290 4876 3292
rect 4630 3238 4632 3290
rect 4812 3238 4814 3290
rect 4568 3236 4574 3238
rect 4630 3236 4654 3238
rect 4710 3236 4734 3238
rect 4790 3236 4814 3238
rect 4870 3236 4876 3238
rect 4568 3216 4876 3236
rect 1854 2748 2162 2768
rect 1854 2746 1860 2748
rect 1916 2746 1940 2748
rect 1996 2746 2020 2748
rect 2076 2746 2100 2748
rect 2156 2746 2162 2748
rect 1916 2694 1918 2746
rect 2098 2694 2100 2746
rect 1854 2692 1860 2694
rect 1916 2692 1940 2694
rect 1996 2692 2020 2694
rect 2076 2692 2100 2694
rect 2156 2692 2162 2694
rect 1854 2672 2162 2692
rect 3664 2748 3972 2768
rect 3664 2746 3670 2748
rect 3726 2746 3750 2748
rect 3806 2746 3830 2748
rect 3886 2746 3910 2748
rect 3966 2746 3972 2748
rect 3726 2694 3728 2746
rect 3908 2694 3910 2746
rect 3664 2692 3670 2694
rect 3726 2692 3750 2694
rect 3806 2692 3830 2694
rect 3886 2692 3910 2694
rect 3966 2692 3972 2694
rect 3664 2672 3972 2692
rect 5473 2748 5781 2768
rect 5473 2746 5479 2748
rect 5535 2746 5559 2748
rect 5615 2746 5639 2748
rect 5695 2746 5719 2748
rect 5775 2746 5781 2748
rect 5535 2694 5537 2746
rect 5717 2694 5719 2746
rect 5473 2692 5479 2694
rect 5535 2692 5559 2694
rect 5615 2692 5639 2694
rect 5695 2692 5719 2694
rect 5775 2692 5781 2694
rect 5473 2672 5781 2692
rect 2759 2204 3067 2224
rect 2759 2202 2765 2204
rect 2821 2202 2845 2204
rect 2901 2202 2925 2204
rect 2981 2202 3005 2204
rect 3061 2202 3067 2204
rect 2821 2150 2823 2202
rect 3003 2150 3005 2202
rect 2759 2148 2765 2150
rect 2821 2148 2845 2150
rect 2901 2148 2925 2150
rect 2981 2148 3005 2150
rect 3061 2148 3067 2150
rect 2759 2128 3067 2148
rect 4568 2204 4876 2224
rect 4568 2202 4574 2204
rect 4630 2202 4654 2204
rect 4710 2202 4734 2204
rect 4790 2202 4814 2204
rect 4870 2202 4876 2204
rect 4630 2150 4632 2202
rect 4812 2150 4814 2202
rect 4568 2148 4574 2150
rect 4630 2148 4654 2150
rect 4710 2148 4734 2150
rect 4790 2148 4814 2150
rect 4870 2148 4876 2150
rect 4568 2128 4876 2148
rect 938 0 994 800
rect 2870 0 2926 800
rect 4802 0 4858 800
rect 6734 0 6790 800
<< via2 >>
rect 2765 7642 2821 7644
rect 2845 7642 2901 7644
rect 2925 7642 2981 7644
rect 3005 7642 3061 7644
rect 2765 7590 2811 7642
rect 2811 7590 2821 7642
rect 2845 7590 2875 7642
rect 2875 7590 2887 7642
rect 2887 7590 2901 7642
rect 2925 7590 2939 7642
rect 2939 7590 2951 7642
rect 2951 7590 2981 7642
rect 3005 7590 3015 7642
rect 3015 7590 3061 7642
rect 2765 7588 2821 7590
rect 2845 7588 2901 7590
rect 2925 7588 2981 7590
rect 3005 7588 3061 7590
rect 4574 7642 4630 7644
rect 4654 7642 4710 7644
rect 4734 7642 4790 7644
rect 4814 7642 4870 7644
rect 4574 7590 4620 7642
rect 4620 7590 4630 7642
rect 4654 7590 4684 7642
rect 4684 7590 4696 7642
rect 4696 7590 4710 7642
rect 4734 7590 4748 7642
rect 4748 7590 4760 7642
rect 4760 7590 4790 7642
rect 4814 7590 4824 7642
rect 4824 7590 4870 7642
rect 4574 7588 4630 7590
rect 4654 7588 4710 7590
rect 4734 7588 4790 7590
rect 4814 7588 4870 7590
rect 1860 7098 1916 7100
rect 1940 7098 1996 7100
rect 2020 7098 2076 7100
rect 2100 7098 2156 7100
rect 1860 7046 1906 7098
rect 1906 7046 1916 7098
rect 1940 7046 1970 7098
rect 1970 7046 1982 7098
rect 1982 7046 1996 7098
rect 2020 7046 2034 7098
rect 2034 7046 2046 7098
rect 2046 7046 2076 7098
rect 2100 7046 2110 7098
rect 2110 7046 2156 7098
rect 1860 7044 1916 7046
rect 1940 7044 1996 7046
rect 2020 7044 2076 7046
rect 2100 7044 2156 7046
rect 3670 7098 3726 7100
rect 3750 7098 3806 7100
rect 3830 7098 3886 7100
rect 3910 7098 3966 7100
rect 3670 7046 3716 7098
rect 3716 7046 3726 7098
rect 3750 7046 3780 7098
rect 3780 7046 3792 7098
rect 3792 7046 3806 7098
rect 3830 7046 3844 7098
rect 3844 7046 3856 7098
rect 3856 7046 3886 7098
rect 3910 7046 3920 7098
rect 3920 7046 3966 7098
rect 3670 7044 3726 7046
rect 3750 7044 3806 7046
rect 3830 7044 3886 7046
rect 3910 7044 3966 7046
rect 5479 7098 5535 7100
rect 5559 7098 5615 7100
rect 5639 7098 5695 7100
rect 5719 7098 5775 7100
rect 5479 7046 5525 7098
rect 5525 7046 5535 7098
rect 5559 7046 5589 7098
rect 5589 7046 5601 7098
rect 5601 7046 5615 7098
rect 5639 7046 5653 7098
rect 5653 7046 5665 7098
rect 5665 7046 5695 7098
rect 5719 7046 5729 7098
rect 5729 7046 5775 7098
rect 5479 7044 5535 7046
rect 5559 7044 5615 7046
rect 5639 7044 5695 7046
rect 5719 7044 5775 7046
rect 2765 6554 2821 6556
rect 2845 6554 2901 6556
rect 2925 6554 2981 6556
rect 3005 6554 3061 6556
rect 2765 6502 2811 6554
rect 2811 6502 2821 6554
rect 2845 6502 2875 6554
rect 2875 6502 2887 6554
rect 2887 6502 2901 6554
rect 2925 6502 2939 6554
rect 2939 6502 2951 6554
rect 2951 6502 2981 6554
rect 3005 6502 3015 6554
rect 3015 6502 3061 6554
rect 2765 6500 2821 6502
rect 2845 6500 2901 6502
rect 2925 6500 2981 6502
rect 3005 6500 3061 6502
rect 4574 6554 4630 6556
rect 4654 6554 4710 6556
rect 4734 6554 4790 6556
rect 4814 6554 4870 6556
rect 4574 6502 4620 6554
rect 4620 6502 4630 6554
rect 4654 6502 4684 6554
rect 4684 6502 4696 6554
rect 4696 6502 4710 6554
rect 4734 6502 4748 6554
rect 4748 6502 4760 6554
rect 4760 6502 4790 6554
rect 4814 6502 4824 6554
rect 4824 6502 4870 6554
rect 4574 6500 4630 6502
rect 4654 6500 4710 6502
rect 4734 6500 4790 6502
rect 4814 6500 4870 6502
rect 1860 6010 1916 6012
rect 1940 6010 1996 6012
rect 2020 6010 2076 6012
rect 2100 6010 2156 6012
rect 1860 5958 1906 6010
rect 1906 5958 1916 6010
rect 1940 5958 1970 6010
rect 1970 5958 1982 6010
rect 1982 5958 1996 6010
rect 2020 5958 2034 6010
rect 2034 5958 2046 6010
rect 2046 5958 2076 6010
rect 2100 5958 2110 6010
rect 2110 5958 2156 6010
rect 1860 5956 1916 5958
rect 1940 5956 1996 5958
rect 2020 5956 2076 5958
rect 2100 5956 2156 5958
rect 3670 6010 3726 6012
rect 3750 6010 3806 6012
rect 3830 6010 3886 6012
rect 3910 6010 3966 6012
rect 3670 5958 3716 6010
rect 3716 5958 3726 6010
rect 3750 5958 3780 6010
rect 3780 5958 3792 6010
rect 3792 5958 3806 6010
rect 3830 5958 3844 6010
rect 3844 5958 3856 6010
rect 3856 5958 3886 6010
rect 3910 5958 3920 6010
rect 3920 5958 3966 6010
rect 3670 5956 3726 5958
rect 3750 5956 3806 5958
rect 3830 5956 3886 5958
rect 3910 5956 3966 5958
rect 5479 6010 5535 6012
rect 5559 6010 5615 6012
rect 5639 6010 5695 6012
rect 5719 6010 5775 6012
rect 5479 5958 5525 6010
rect 5525 5958 5535 6010
rect 5559 5958 5589 6010
rect 5589 5958 5601 6010
rect 5601 5958 5615 6010
rect 5639 5958 5653 6010
rect 5653 5958 5665 6010
rect 5665 5958 5695 6010
rect 5719 5958 5729 6010
rect 5729 5958 5775 6010
rect 5479 5956 5535 5958
rect 5559 5956 5615 5958
rect 5639 5956 5695 5958
rect 5719 5956 5775 5958
rect 2765 5466 2821 5468
rect 2845 5466 2901 5468
rect 2925 5466 2981 5468
rect 3005 5466 3061 5468
rect 2765 5414 2811 5466
rect 2811 5414 2821 5466
rect 2845 5414 2875 5466
rect 2875 5414 2887 5466
rect 2887 5414 2901 5466
rect 2925 5414 2939 5466
rect 2939 5414 2951 5466
rect 2951 5414 2981 5466
rect 3005 5414 3015 5466
rect 3015 5414 3061 5466
rect 2765 5412 2821 5414
rect 2845 5412 2901 5414
rect 2925 5412 2981 5414
rect 3005 5412 3061 5414
rect 4574 5466 4630 5468
rect 4654 5466 4710 5468
rect 4734 5466 4790 5468
rect 4814 5466 4870 5468
rect 4574 5414 4620 5466
rect 4620 5414 4630 5466
rect 4654 5414 4684 5466
rect 4684 5414 4696 5466
rect 4696 5414 4710 5466
rect 4734 5414 4748 5466
rect 4748 5414 4760 5466
rect 4760 5414 4790 5466
rect 4814 5414 4824 5466
rect 4824 5414 4870 5466
rect 4574 5412 4630 5414
rect 4654 5412 4710 5414
rect 4734 5412 4790 5414
rect 4814 5412 4870 5414
rect 5906 4972 5908 4992
rect 5908 4972 5960 4992
rect 5960 4972 5962 4992
rect 1860 4922 1916 4924
rect 1940 4922 1996 4924
rect 2020 4922 2076 4924
rect 2100 4922 2156 4924
rect 1860 4870 1906 4922
rect 1906 4870 1916 4922
rect 1940 4870 1970 4922
rect 1970 4870 1982 4922
rect 1982 4870 1996 4922
rect 2020 4870 2034 4922
rect 2034 4870 2046 4922
rect 2046 4870 2076 4922
rect 2100 4870 2110 4922
rect 2110 4870 2156 4922
rect 1860 4868 1916 4870
rect 1940 4868 1996 4870
rect 2020 4868 2076 4870
rect 2100 4868 2156 4870
rect 3670 4922 3726 4924
rect 3750 4922 3806 4924
rect 3830 4922 3886 4924
rect 3910 4922 3966 4924
rect 3670 4870 3716 4922
rect 3716 4870 3726 4922
rect 3750 4870 3780 4922
rect 3780 4870 3792 4922
rect 3792 4870 3806 4922
rect 3830 4870 3844 4922
rect 3844 4870 3856 4922
rect 3856 4870 3886 4922
rect 3910 4870 3920 4922
rect 3920 4870 3966 4922
rect 3670 4868 3726 4870
rect 3750 4868 3806 4870
rect 3830 4868 3886 4870
rect 3910 4868 3966 4870
rect 5906 4936 5962 4972
rect 5479 4922 5535 4924
rect 5559 4922 5615 4924
rect 5639 4922 5695 4924
rect 5719 4922 5775 4924
rect 5479 4870 5525 4922
rect 5525 4870 5535 4922
rect 5559 4870 5589 4922
rect 5589 4870 5601 4922
rect 5601 4870 5615 4922
rect 5639 4870 5653 4922
rect 5653 4870 5665 4922
rect 5665 4870 5695 4922
rect 5719 4870 5729 4922
rect 5729 4870 5775 4922
rect 5479 4868 5535 4870
rect 5559 4868 5615 4870
rect 5639 4868 5695 4870
rect 5719 4868 5775 4870
rect 2765 4378 2821 4380
rect 2845 4378 2901 4380
rect 2925 4378 2981 4380
rect 3005 4378 3061 4380
rect 2765 4326 2811 4378
rect 2811 4326 2821 4378
rect 2845 4326 2875 4378
rect 2875 4326 2887 4378
rect 2887 4326 2901 4378
rect 2925 4326 2939 4378
rect 2939 4326 2951 4378
rect 2951 4326 2981 4378
rect 3005 4326 3015 4378
rect 3015 4326 3061 4378
rect 2765 4324 2821 4326
rect 2845 4324 2901 4326
rect 2925 4324 2981 4326
rect 3005 4324 3061 4326
rect 4574 4378 4630 4380
rect 4654 4378 4710 4380
rect 4734 4378 4790 4380
rect 4814 4378 4870 4380
rect 4574 4326 4620 4378
rect 4620 4326 4630 4378
rect 4654 4326 4684 4378
rect 4684 4326 4696 4378
rect 4696 4326 4710 4378
rect 4734 4326 4748 4378
rect 4748 4326 4760 4378
rect 4760 4326 4790 4378
rect 4814 4326 4824 4378
rect 4824 4326 4870 4378
rect 4574 4324 4630 4326
rect 4654 4324 4710 4326
rect 4734 4324 4790 4326
rect 4814 4324 4870 4326
rect 1860 3834 1916 3836
rect 1940 3834 1996 3836
rect 2020 3834 2076 3836
rect 2100 3834 2156 3836
rect 1860 3782 1906 3834
rect 1906 3782 1916 3834
rect 1940 3782 1970 3834
rect 1970 3782 1982 3834
rect 1982 3782 1996 3834
rect 2020 3782 2034 3834
rect 2034 3782 2046 3834
rect 2046 3782 2076 3834
rect 2100 3782 2110 3834
rect 2110 3782 2156 3834
rect 1860 3780 1916 3782
rect 1940 3780 1996 3782
rect 2020 3780 2076 3782
rect 2100 3780 2156 3782
rect 3670 3834 3726 3836
rect 3750 3834 3806 3836
rect 3830 3834 3886 3836
rect 3910 3834 3966 3836
rect 3670 3782 3716 3834
rect 3716 3782 3726 3834
rect 3750 3782 3780 3834
rect 3780 3782 3792 3834
rect 3792 3782 3806 3834
rect 3830 3782 3844 3834
rect 3844 3782 3856 3834
rect 3856 3782 3886 3834
rect 3910 3782 3920 3834
rect 3920 3782 3966 3834
rect 3670 3780 3726 3782
rect 3750 3780 3806 3782
rect 3830 3780 3886 3782
rect 3910 3780 3966 3782
rect 5479 3834 5535 3836
rect 5559 3834 5615 3836
rect 5639 3834 5695 3836
rect 5719 3834 5775 3836
rect 5479 3782 5525 3834
rect 5525 3782 5535 3834
rect 5559 3782 5589 3834
rect 5589 3782 5601 3834
rect 5601 3782 5615 3834
rect 5639 3782 5653 3834
rect 5653 3782 5665 3834
rect 5665 3782 5695 3834
rect 5719 3782 5729 3834
rect 5729 3782 5775 3834
rect 5479 3780 5535 3782
rect 5559 3780 5615 3782
rect 5639 3780 5695 3782
rect 5719 3780 5775 3782
rect 2765 3290 2821 3292
rect 2845 3290 2901 3292
rect 2925 3290 2981 3292
rect 3005 3290 3061 3292
rect 2765 3238 2811 3290
rect 2811 3238 2821 3290
rect 2845 3238 2875 3290
rect 2875 3238 2887 3290
rect 2887 3238 2901 3290
rect 2925 3238 2939 3290
rect 2939 3238 2951 3290
rect 2951 3238 2981 3290
rect 3005 3238 3015 3290
rect 3015 3238 3061 3290
rect 2765 3236 2821 3238
rect 2845 3236 2901 3238
rect 2925 3236 2981 3238
rect 3005 3236 3061 3238
rect 4574 3290 4630 3292
rect 4654 3290 4710 3292
rect 4734 3290 4790 3292
rect 4814 3290 4870 3292
rect 4574 3238 4620 3290
rect 4620 3238 4630 3290
rect 4654 3238 4684 3290
rect 4684 3238 4696 3290
rect 4696 3238 4710 3290
rect 4734 3238 4748 3290
rect 4748 3238 4760 3290
rect 4760 3238 4790 3290
rect 4814 3238 4824 3290
rect 4824 3238 4870 3290
rect 4574 3236 4630 3238
rect 4654 3236 4710 3238
rect 4734 3236 4790 3238
rect 4814 3236 4870 3238
rect 1860 2746 1916 2748
rect 1940 2746 1996 2748
rect 2020 2746 2076 2748
rect 2100 2746 2156 2748
rect 1860 2694 1906 2746
rect 1906 2694 1916 2746
rect 1940 2694 1970 2746
rect 1970 2694 1982 2746
rect 1982 2694 1996 2746
rect 2020 2694 2034 2746
rect 2034 2694 2046 2746
rect 2046 2694 2076 2746
rect 2100 2694 2110 2746
rect 2110 2694 2156 2746
rect 1860 2692 1916 2694
rect 1940 2692 1996 2694
rect 2020 2692 2076 2694
rect 2100 2692 2156 2694
rect 3670 2746 3726 2748
rect 3750 2746 3806 2748
rect 3830 2746 3886 2748
rect 3910 2746 3966 2748
rect 3670 2694 3716 2746
rect 3716 2694 3726 2746
rect 3750 2694 3780 2746
rect 3780 2694 3792 2746
rect 3792 2694 3806 2746
rect 3830 2694 3844 2746
rect 3844 2694 3856 2746
rect 3856 2694 3886 2746
rect 3910 2694 3920 2746
rect 3920 2694 3966 2746
rect 3670 2692 3726 2694
rect 3750 2692 3806 2694
rect 3830 2692 3886 2694
rect 3910 2692 3966 2694
rect 5479 2746 5535 2748
rect 5559 2746 5615 2748
rect 5639 2746 5695 2748
rect 5719 2746 5775 2748
rect 5479 2694 5525 2746
rect 5525 2694 5535 2746
rect 5559 2694 5589 2746
rect 5589 2694 5601 2746
rect 5601 2694 5615 2746
rect 5639 2694 5653 2746
rect 5653 2694 5665 2746
rect 5665 2694 5695 2746
rect 5719 2694 5729 2746
rect 5729 2694 5775 2746
rect 5479 2692 5535 2694
rect 5559 2692 5615 2694
rect 5639 2692 5695 2694
rect 5719 2692 5775 2694
rect 2765 2202 2821 2204
rect 2845 2202 2901 2204
rect 2925 2202 2981 2204
rect 3005 2202 3061 2204
rect 2765 2150 2811 2202
rect 2811 2150 2821 2202
rect 2845 2150 2875 2202
rect 2875 2150 2887 2202
rect 2887 2150 2901 2202
rect 2925 2150 2939 2202
rect 2939 2150 2951 2202
rect 2951 2150 2981 2202
rect 3005 2150 3015 2202
rect 3015 2150 3061 2202
rect 2765 2148 2821 2150
rect 2845 2148 2901 2150
rect 2925 2148 2981 2150
rect 3005 2148 3061 2150
rect 4574 2202 4630 2204
rect 4654 2202 4710 2204
rect 4734 2202 4790 2204
rect 4814 2202 4870 2204
rect 4574 2150 4620 2202
rect 4620 2150 4630 2202
rect 4654 2150 4684 2202
rect 4684 2150 4696 2202
rect 4696 2150 4710 2202
rect 4734 2150 4748 2202
rect 4748 2150 4760 2202
rect 4760 2150 4790 2202
rect 4814 2150 4824 2202
rect 4824 2150 4870 2202
rect 4574 2148 4630 2150
rect 4654 2148 4710 2150
rect 4734 2148 4790 2150
rect 4814 2148 4870 2150
<< metal3 >>
rect 6888 8168 7688 8288
rect 2753 7648 3073 7649
rect 2753 7584 2761 7648
rect 2825 7584 2841 7648
rect 2905 7584 2921 7648
rect 2985 7584 3001 7648
rect 3065 7584 3073 7648
rect 2753 7583 3073 7584
rect 4562 7648 4882 7649
rect 4562 7584 4570 7648
rect 4634 7584 4650 7648
rect 4714 7584 4730 7648
rect 4794 7584 4810 7648
rect 4874 7584 4882 7648
rect 4562 7583 4882 7584
rect 0 7352 800 7472
rect 1848 7104 2168 7105
rect 1848 7040 1856 7104
rect 1920 7040 1936 7104
rect 2000 7040 2016 7104
rect 2080 7040 2096 7104
rect 2160 7040 2168 7104
rect 1848 7039 2168 7040
rect 3658 7104 3978 7105
rect 3658 7040 3666 7104
rect 3730 7040 3746 7104
rect 3810 7040 3826 7104
rect 3890 7040 3906 7104
rect 3970 7040 3978 7104
rect 3658 7039 3978 7040
rect 5467 7104 5787 7105
rect 5467 7040 5475 7104
rect 5539 7040 5555 7104
rect 5619 7040 5635 7104
rect 5699 7040 5715 7104
rect 5779 7040 5787 7104
rect 5467 7039 5787 7040
rect 2753 6560 3073 6561
rect 2753 6496 2761 6560
rect 2825 6496 2841 6560
rect 2905 6496 2921 6560
rect 2985 6496 3001 6560
rect 3065 6496 3073 6560
rect 2753 6495 3073 6496
rect 4562 6560 4882 6561
rect 4562 6496 4570 6560
rect 4634 6496 4650 6560
rect 4714 6496 4730 6560
rect 4794 6496 4810 6560
rect 4874 6496 4882 6560
rect 4562 6495 4882 6496
rect 1848 6016 2168 6017
rect 1848 5952 1856 6016
rect 1920 5952 1936 6016
rect 2000 5952 2016 6016
rect 2080 5952 2096 6016
rect 2160 5952 2168 6016
rect 1848 5951 2168 5952
rect 3658 6016 3978 6017
rect 3658 5952 3666 6016
rect 3730 5952 3746 6016
rect 3810 5952 3826 6016
rect 3890 5952 3906 6016
rect 3970 5952 3978 6016
rect 3658 5951 3978 5952
rect 5467 6016 5787 6017
rect 5467 5952 5475 6016
rect 5539 5952 5555 6016
rect 5619 5952 5635 6016
rect 5699 5952 5715 6016
rect 5779 5952 5787 6016
rect 5467 5951 5787 5952
rect 2753 5472 3073 5473
rect 2753 5408 2761 5472
rect 2825 5408 2841 5472
rect 2905 5408 2921 5472
rect 2985 5408 3001 5472
rect 3065 5408 3073 5472
rect 2753 5407 3073 5408
rect 4562 5472 4882 5473
rect 4562 5408 4570 5472
rect 4634 5408 4650 5472
rect 4714 5408 4730 5472
rect 4794 5408 4810 5472
rect 4874 5408 4882 5472
rect 4562 5407 4882 5408
rect 5901 4994 5967 4997
rect 6888 4994 7688 5024
rect 5901 4992 7688 4994
rect 5901 4936 5906 4992
rect 5962 4936 7688 4992
rect 5901 4934 7688 4936
rect 5901 4931 5967 4934
rect 1848 4928 2168 4929
rect 1848 4864 1856 4928
rect 1920 4864 1936 4928
rect 2000 4864 2016 4928
rect 2080 4864 2096 4928
rect 2160 4864 2168 4928
rect 1848 4863 2168 4864
rect 3658 4928 3978 4929
rect 3658 4864 3666 4928
rect 3730 4864 3746 4928
rect 3810 4864 3826 4928
rect 3890 4864 3906 4928
rect 3970 4864 3978 4928
rect 3658 4863 3978 4864
rect 5467 4928 5787 4929
rect 5467 4864 5475 4928
rect 5539 4864 5555 4928
rect 5619 4864 5635 4928
rect 5699 4864 5715 4928
rect 5779 4864 5787 4928
rect 6888 4904 7688 4934
rect 5467 4863 5787 4864
rect 2753 4384 3073 4385
rect 2753 4320 2761 4384
rect 2825 4320 2841 4384
rect 2905 4320 2921 4384
rect 2985 4320 3001 4384
rect 3065 4320 3073 4384
rect 2753 4319 3073 4320
rect 4562 4384 4882 4385
rect 4562 4320 4570 4384
rect 4634 4320 4650 4384
rect 4714 4320 4730 4384
rect 4794 4320 4810 4384
rect 4874 4320 4882 4384
rect 4562 4319 4882 4320
rect 1848 3840 2168 3841
rect 1848 3776 1856 3840
rect 1920 3776 1936 3840
rect 2000 3776 2016 3840
rect 2080 3776 2096 3840
rect 2160 3776 2168 3840
rect 1848 3775 2168 3776
rect 3658 3840 3978 3841
rect 3658 3776 3666 3840
rect 3730 3776 3746 3840
rect 3810 3776 3826 3840
rect 3890 3776 3906 3840
rect 3970 3776 3978 3840
rect 3658 3775 3978 3776
rect 5467 3840 5787 3841
rect 5467 3776 5475 3840
rect 5539 3776 5555 3840
rect 5619 3776 5635 3840
rect 5699 3776 5715 3840
rect 5779 3776 5787 3840
rect 5467 3775 5787 3776
rect 2753 3296 3073 3297
rect 2753 3232 2761 3296
rect 2825 3232 2841 3296
rect 2905 3232 2921 3296
rect 2985 3232 3001 3296
rect 3065 3232 3073 3296
rect 2753 3231 3073 3232
rect 4562 3296 4882 3297
rect 4562 3232 4570 3296
rect 4634 3232 4650 3296
rect 4714 3232 4730 3296
rect 4794 3232 4810 3296
rect 4874 3232 4882 3296
rect 4562 3231 4882 3232
rect 1848 2752 2168 2753
rect 1848 2688 1856 2752
rect 1920 2688 1936 2752
rect 2000 2688 2016 2752
rect 2080 2688 2096 2752
rect 2160 2688 2168 2752
rect 1848 2687 2168 2688
rect 3658 2752 3978 2753
rect 3658 2688 3666 2752
rect 3730 2688 3746 2752
rect 3810 2688 3826 2752
rect 3890 2688 3906 2752
rect 3970 2688 3978 2752
rect 3658 2687 3978 2688
rect 5467 2752 5787 2753
rect 5467 2688 5475 2752
rect 5539 2688 5555 2752
rect 5619 2688 5635 2752
rect 5699 2688 5715 2752
rect 5779 2688 5787 2752
rect 5467 2687 5787 2688
rect 0 2456 800 2576
rect 2753 2208 3073 2209
rect 2753 2144 2761 2208
rect 2825 2144 2841 2208
rect 2905 2144 2921 2208
rect 2985 2144 3001 2208
rect 3065 2144 3073 2208
rect 2753 2143 3073 2144
rect 4562 2208 4882 2209
rect 4562 2144 4570 2208
rect 4634 2144 4650 2208
rect 4714 2144 4730 2208
rect 4794 2144 4810 2208
rect 4874 2144 4882 2208
rect 4562 2143 4882 2144
rect 6888 1640 7688 1760
<< via3 >>
rect 2761 7644 2825 7648
rect 2761 7588 2765 7644
rect 2765 7588 2821 7644
rect 2821 7588 2825 7644
rect 2761 7584 2825 7588
rect 2841 7644 2905 7648
rect 2841 7588 2845 7644
rect 2845 7588 2901 7644
rect 2901 7588 2905 7644
rect 2841 7584 2905 7588
rect 2921 7644 2985 7648
rect 2921 7588 2925 7644
rect 2925 7588 2981 7644
rect 2981 7588 2985 7644
rect 2921 7584 2985 7588
rect 3001 7644 3065 7648
rect 3001 7588 3005 7644
rect 3005 7588 3061 7644
rect 3061 7588 3065 7644
rect 3001 7584 3065 7588
rect 4570 7644 4634 7648
rect 4570 7588 4574 7644
rect 4574 7588 4630 7644
rect 4630 7588 4634 7644
rect 4570 7584 4634 7588
rect 4650 7644 4714 7648
rect 4650 7588 4654 7644
rect 4654 7588 4710 7644
rect 4710 7588 4714 7644
rect 4650 7584 4714 7588
rect 4730 7644 4794 7648
rect 4730 7588 4734 7644
rect 4734 7588 4790 7644
rect 4790 7588 4794 7644
rect 4730 7584 4794 7588
rect 4810 7644 4874 7648
rect 4810 7588 4814 7644
rect 4814 7588 4870 7644
rect 4870 7588 4874 7644
rect 4810 7584 4874 7588
rect 1856 7100 1920 7104
rect 1856 7044 1860 7100
rect 1860 7044 1916 7100
rect 1916 7044 1920 7100
rect 1856 7040 1920 7044
rect 1936 7100 2000 7104
rect 1936 7044 1940 7100
rect 1940 7044 1996 7100
rect 1996 7044 2000 7100
rect 1936 7040 2000 7044
rect 2016 7100 2080 7104
rect 2016 7044 2020 7100
rect 2020 7044 2076 7100
rect 2076 7044 2080 7100
rect 2016 7040 2080 7044
rect 2096 7100 2160 7104
rect 2096 7044 2100 7100
rect 2100 7044 2156 7100
rect 2156 7044 2160 7100
rect 2096 7040 2160 7044
rect 3666 7100 3730 7104
rect 3666 7044 3670 7100
rect 3670 7044 3726 7100
rect 3726 7044 3730 7100
rect 3666 7040 3730 7044
rect 3746 7100 3810 7104
rect 3746 7044 3750 7100
rect 3750 7044 3806 7100
rect 3806 7044 3810 7100
rect 3746 7040 3810 7044
rect 3826 7100 3890 7104
rect 3826 7044 3830 7100
rect 3830 7044 3886 7100
rect 3886 7044 3890 7100
rect 3826 7040 3890 7044
rect 3906 7100 3970 7104
rect 3906 7044 3910 7100
rect 3910 7044 3966 7100
rect 3966 7044 3970 7100
rect 3906 7040 3970 7044
rect 5475 7100 5539 7104
rect 5475 7044 5479 7100
rect 5479 7044 5535 7100
rect 5535 7044 5539 7100
rect 5475 7040 5539 7044
rect 5555 7100 5619 7104
rect 5555 7044 5559 7100
rect 5559 7044 5615 7100
rect 5615 7044 5619 7100
rect 5555 7040 5619 7044
rect 5635 7100 5699 7104
rect 5635 7044 5639 7100
rect 5639 7044 5695 7100
rect 5695 7044 5699 7100
rect 5635 7040 5699 7044
rect 5715 7100 5779 7104
rect 5715 7044 5719 7100
rect 5719 7044 5775 7100
rect 5775 7044 5779 7100
rect 5715 7040 5779 7044
rect 2761 6556 2825 6560
rect 2761 6500 2765 6556
rect 2765 6500 2821 6556
rect 2821 6500 2825 6556
rect 2761 6496 2825 6500
rect 2841 6556 2905 6560
rect 2841 6500 2845 6556
rect 2845 6500 2901 6556
rect 2901 6500 2905 6556
rect 2841 6496 2905 6500
rect 2921 6556 2985 6560
rect 2921 6500 2925 6556
rect 2925 6500 2981 6556
rect 2981 6500 2985 6556
rect 2921 6496 2985 6500
rect 3001 6556 3065 6560
rect 3001 6500 3005 6556
rect 3005 6500 3061 6556
rect 3061 6500 3065 6556
rect 3001 6496 3065 6500
rect 4570 6556 4634 6560
rect 4570 6500 4574 6556
rect 4574 6500 4630 6556
rect 4630 6500 4634 6556
rect 4570 6496 4634 6500
rect 4650 6556 4714 6560
rect 4650 6500 4654 6556
rect 4654 6500 4710 6556
rect 4710 6500 4714 6556
rect 4650 6496 4714 6500
rect 4730 6556 4794 6560
rect 4730 6500 4734 6556
rect 4734 6500 4790 6556
rect 4790 6500 4794 6556
rect 4730 6496 4794 6500
rect 4810 6556 4874 6560
rect 4810 6500 4814 6556
rect 4814 6500 4870 6556
rect 4870 6500 4874 6556
rect 4810 6496 4874 6500
rect 1856 6012 1920 6016
rect 1856 5956 1860 6012
rect 1860 5956 1916 6012
rect 1916 5956 1920 6012
rect 1856 5952 1920 5956
rect 1936 6012 2000 6016
rect 1936 5956 1940 6012
rect 1940 5956 1996 6012
rect 1996 5956 2000 6012
rect 1936 5952 2000 5956
rect 2016 6012 2080 6016
rect 2016 5956 2020 6012
rect 2020 5956 2076 6012
rect 2076 5956 2080 6012
rect 2016 5952 2080 5956
rect 2096 6012 2160 6016
rect 2096 5956 2100 6012
rect 2100 5956 2156 6012
rect 2156 5956 2160 6012
rect 2096 5952 2160 5956
rect 3666 6012 3730 6016
rect 3666 5956 3670 6012
rect 3670 5956 3726 6012
rect 3726 5956 3730 6012
rect 3666 5952 3730 5956
rect 3746 6012 3810 6016
rect 3746 5956 3750 6012
rect 3750 5956 3806 6012
rect 3806 5956 3810 6012
rect 3746 5952 3810 5956
rect 3826 6012 3890 6016
rect 3826 5956 3830 6012
rect 3830 5956 3886 6012
rect 3886 5956 3890 6012
rect 3826 5952 3890 5956
rect 3906 6012 3970 6016
rect 3906 5956 3910 6012
rect 3910 5956 3966 6012
rect 3966 5956 3970 6012
rect 3906 5952 3970 5956
rect 5475 6012 5539 6016
rect 5475 5956 5479 6012
rect 5479 5956 5535 6012
rect 5535 5956 5539 6012
rect 5475 5952 5539 5956
rect 5555 6012 5619 6016
rect 5555 5956 5559 6012
rect 5559 5956 5615 6012
rect 5615 5956 5619 6012
rect 5555 5952 5619 5956
rect 5635 6012 5699 6016
rect 5635 5956 5639 6012
rect 5639 5956 5695 6012
rect 5695 5956 5699 6012
rect 5635 5952 5699 5956
rect 5715 6012 5779 6016
rect 5715 5956 5719 6012
rect 5719 5956 5775 6012
rect 5775 5956 5779 6012
rect 5715 5952 5779 5956
rect 2761 5468 2825 5472
rect 2761 5412 2765 5468
rect 2765 5412 2821 5468
rect 2821 5412 2825 5468
rect 2761 5408 2825 5412
rect 2841 5468 2905 5472
rect 2841 5412 2845 5468
rect 2845 5412 2901 5468
rect 2901 5412 2905 5468
rect 2841 5408 2905 5412
rect 2921 5468 2985 5472
rect 2921 5412 2925 5468
rect 2925 5412 2981 5468
rect 2981 5412 2985 5468
rect 2921 5408 2985 5412
rect 3001 5468 3065 5472
rect 3001 5412 3005 5468
rect 3005 5412 3061 5468
rect 3061 5412 3065 5468
rect 3001 5408 3065 5412
rect 4570 5468 4634 5472
rect 4570 5412 4574 5468
rect 4574 5412 4630 5468
rect 4630 5412 4634 5468
rect 4570 5408 4634 5412
rect 4650 5468 4714 5472
rect 4650 5412 4654 5468
rect 4654 5412 4710 5468
rect 4710 5412 4714 5468
rect 4650 5408 4714 5412
rect 4730 5468 4794 5472
rect 4730 5412 4734 5468
rect 4734 5412 4790 5468
rect 4790 5412 4794 5468
rect 4730 5408 4794 5412
rect 4810 5468 4874 5472
rect 4810 5412 4814 5468
rect 4814 5412 4870 5468
rect 4870 5412 4874 5468
rect 4810 5408 4874 5412
rect 1856 4924 1920 4928
rect 1856 4868 1860 4924
rect 1860 4868 1916 4924
rect 1916 4868 1920 4924
rect 1856 4864 1920 4868
rect 1936 4924 2000 4928
rect 1936 4868 1940 4924
rect 1940 4868 1996 4924
rect 1996 4868 2000 4924
rect 1936 4864 2000 4868
rect 2016 4924 2080 4928
rect 2016 4868 2020 4924
rect 2020 4868 2076 4924
rect 2076 4868 2080 4924
rect 2016 4864 2080 4868
rect 2096 4924 2160 4928
rect 2096 4868 2100 4924
rect 2100 4868 2156 4924
rect 2156 4868 2160 4924
rect 2096 4864 2160 4868
rect 3666 4924 3730 4928
rect 3666 4868 3670 4924
rect 3670 4868 3726 4924
rect 3726 4868 3730 4924
rect 3666 4864 3730 4868
rect 3746 4924 3810 4928
rect 3746 4868 3750 4924
rect 3750 4868 3806 4924
rect 3806 4868 3810 4924
rect 3746 4864 3810 4868
rect 3826 4924 3890 4928
rect 3826 4868 3830 4924
rect 3830 4868 3886 4924
rect 3886 4868 3890 4924
rect 3826 4864 3890 4868
rect 3906 4924 3970 4928
rect 3906 4868 3910 4924
rect 3910 4868 3966 4924
rect 3966 4868 3970 4924
rect 3906 4864 3970 4868
rect 5475 4924 5539 4928
rect 5475 4868 5479 4924
rect 5479 4868 5535 4924
rect 5535 4868 5539 4924
rect 5475 4864 5539 4868
rect 5555 4924 5619 4928
rect 5555 4868 5559 4924
rect 5559 4868 5615 4924
rect 5615 4868 5619 4924
rect 5555 4864 5619 4868
rect 5635 4924 5699 4928
rect 5635 4868 5639 4924
rect 5639 4868 5695 4924
rect 5695 4868 5699 4924
rect 5635 4864 5699 4868
rect 5715 4924 5779 4928
rect 5715 4868 5719 4924
rect 5719 4868 5775 4924
rect 5775 4868 5779 4924
rect 5715 4864 5779 4868
rect 2761 4380 2825 4384
rect 2761 4324 2765 4380
rect 2765 4324 2821 4380
rect 2821 4324 2825 4380
rect 2761 4320 2825 4324
rect 2841 4380 2905 4384
rect 2841 4324 2845 4380
rect 2845 4324 2901 4380
rect 2901 4324 2905 4380
rect 2841 4320 2905 4324
rect 2921 4380 2985 4384
rect 2921 4324 2925 4380
rect 2925 4324 2981 4380
rect 2981 4324 2985 4380
rect 2921 4320 2985 4324
rect 3001 4380 3065 4384
rect 3001 4324 3005 4380
rect 3005 4324 3061 4380
rect 3061 4324 3065 4380
rect 3001 4320 3065 4324
rect 4570 4380 4634 4384
rect 4570 4324 4574 4380
rect 4574 4324 4630 4380
rect 4630 4324 4634 4380
rect 4570 4320 4634 4324
rect 4650 4380 4714 4384
rect 4650 4324 4654 4380
rect 4654 4324 4710 4380
rect 4710 4324 4714 4380
rect 4650 4320 4714 4324
rect 4730 4380 4794 4384
rect 4730 4324 4734 4380
rect 4734 4324 4790 4380
rect 4790 4324 4794 4380
rect 4730 4320 4794 4324
rect 4810 4380 4874 4384
rect 4810 4324 4814 4380
rect 4814 4324 4870 4380
rect 4870 4324 4874 4380
rect 4810 4320 4874 4324
rect 1856 3836 1920 3840
rect 1856 3780 1860 3836
rect 1860 3780 1916 3836
rect 1916 3780 1920 3836
rect 1856 3776 1920 3780
rect 1936 3836 2000 3840
rect 1936 3780 1940 3836
rect 1940 3780 1996 3836
rect 1996 3780 2000 3836
rect 1936 3776 2000 3780
rect 2016 3836 2080 3840
rect 2016 3780 2020 3836
rect 2020 3780 2076 3836
rect 2076 3780 2080 3836
rect 2016 3776 2080 3780
rect 2096 3836 2160 3840
rect 2096 3780 2100 3836
rect 2100 3780 2156 3836
rect 2156 3780 2160 3836
rect 2096 3776 2160 3780
rect 3666 3836 3730 3840
rect 3666 3780 3670 3836
rect 3670 3780 3726 3836
rect 3726 3780 3730 3836
rect 3666 3776 3730 3780
rect 3746 3836 3810 3840
rect 3746 3780 3750 3836
rect 3750 3780 3806 3836
rect 3806 3780 3810 3836
rect 3746 3776 3810 3780
rect 3826 3836 3890 3840
rect 3826 3780 3830 3836
rect 3830 3780 3886 3836
rect 3886 3780 3890 3836
rect 3826 3776 3890 3780
rect 3906 3836 3970 3840
rect 3906 3780 3910 3836
rect 3910 3780 3966 3836
rect 3966 3780 3970 3836
rect 3906 3776 3970 3780
rect 5475 3836 5539 3840
rect 5475 3780 5479 3836
rect 5479 3780 5535 3836
rect 5535 3780 5539 3836
rect 5475 3776 5539 3780
rect 5555 3836 5619 3840
rect 5555 3780 5559 3836
rect 5559 3780 5615 3836
rect 5615 3780 5619 3836
rect 5555 3776 5619 3780
rect 5635 3836 5699 3840
rect 5635 3780 5639 3836
rect 5639 3780 5695 3836
rect 5695 3780 5699 3836
rect 5635 3776 5699 3780
rect 5715 3836 5779 3840
rect 5715 3780 5719 3836
rect 5719 3780 5775 3836
rect 5775 3780 5779 3836
rect 5715 3776 5779 3780
rect 2761 3292 2825 3296
rect 2761 3236 2765 3292
rect 2765 3236 2821 3292
rect 2821 3236 2825 3292
rect 2761 3232 2825 3236
rect 2841 3292 2905 3296
rect 2841 3236 2845 3292
rect 2845 3236 2901 3292
rect 2901 3236 2905 3292
rect 2841 3232 2905 3236
rect 2921 3292 2985 3296
rect 2921 3236 2925 3292
rect 2925 3236 2981 3292
rect 2981 3236 2985 3292
rect 2921 3232 2985 3236
rect 3001 3292 3065 3296
rect 3001 3236 3005 3292
rect 3005 3236 3061 3292
rect 3061 3236 3065 3292
rect 3001 3232 3065 3236
rect 4570 3292 4634 3296
rect 4570 3236 4574 3292
rect 4574 3236 4630 3292
rect 4630 3236 4634 3292
rect 4570 3232 4634 3236
rect 4650 3292 4714 3296
rect 4650 3236 4654 3292
rect 4654 3236 4710 3292
rect 4710 3236 4714 3292
rect 4650 3232 4714 3236
rect 4730 3292 4794 3296
rect 4730 3236 4734 3292
rect 4734 3236 4790 3292
rect 4790 3236 4794 3292
rect 4730 3232 4794 3236
rect 4810 3292 4874 3296
rect 4810 3236 4814 3292
rect 4814 3236 4870 3292
rect 4870 3236 4874 3292
rect 4810 3232 4874 3236
rect 1856 2748 1920 2752
rect 1856 2692 1860 2748
rect 1860 2692 1916 2748
rect 1916 2692 1920 2748
rect 1856 2688 1920 2692
rect 1936 2748 2000 2752
rect 1936 2692 1940 2748
rect 1940 2692 1996 2748
rect 1996 2692 2000 2748
rect 1936 2688 2000 2692
rect 2016 2748 2080 2752
rect 2016 2692 2020 2748
rect 2020 2692 2076 2748
rect 2076 2692 2080 2748
rect 2016 2688 2080 2692
rect 2096 2748 2160 2752
rect 2096 2692 2100 2748
rect 2100 2692 2156 2748
rect 2156 2692 2160 2748
rect 2096 2688 2160 2692
rect 3666 2748 3730 2752
rect 3666 2692 3670 2748
rect 3670 2692 3726 2748
rect 3726 2692 3730 2748
rect 3666 2688 3730 2692
rect 3746 2748 3810 2752
rect 3746 2692 3750 2748
rect 3750 2692 3806 2748
rect 3806 2692 3810 2748
rect 3746 2688 3810 2692
rect 3826 2748 3890 2752
rect 3826 2692 3830 2748
rect 3830 2692 3886 2748
rect 3886 2692 3890 2748
rect 3826 2688 3890 2692
rect 3906 2748 3970 2752
rect 3906 2692 3910 2748
rect 3910 2692 3966 2748
rect 3966 2692 3970 2748
rect 3906 2688 3970 2692
rect 5475 2748 5539 2752
rect 5475 2692 5479 2748
rect 5479 2692 5535 2748
rect 5535 2692 5539 2748
rect 5475 2688 5539 2692
rect 5555 2748 5619 2752
rect 5555 2692 5559 2748
rect 5559 2692 5615 2748
rect 5615 2692 5619 2748
rect 5555 2688 5619 2692
rect 5635 2748 5699 2752
rect 5635 2692 5639 2748
rect 5639 2692 5695 2748
rect 5695 2692 5699 2748
rect 5635 2688 5699 2692
rect 5715 2748 5779 2752
rect 5715 2692 5719 2748
rect 5719 2692 5775 2748
rect 5775 2692 5779 2748
rect 5715 2688 5779 2692
rect 2761 2204 2825 2208
rect 2761 2148 2765 2204
rect 2765 2148 2821 2204
rect 2821 2148 2825 2204
rect 2761 2144 2825 2148
rect 2841 2204 2905 2208
rect 2841 2148 2845 2204
rect 2845 2148 2901 2204
rect 2901 2148 2905 2204
rect 2841 2144 2905 2148
rect 2921 2204 2985 2208
rect 2921 2148 2925 2204
rect 2925 2148 2981 2204
rect 2981 2148 2985 2204
rect 2921 2144 2985 2148
rect 3001 2204 3065 2208
rect 3001 2148 3005 2204
rect 3005 2148 3061 2204
rect 3061 2148 3065 2204
rect 3001 2144 3065 2148
rect 4570 2204 4634 2208
rect 4570 2148 4574 2204
rect 4574 2148 4630 2204
rect 4630 2148 4634 2204
rect 4570 2144 4634 2148
rect 4650 2204 4714 2208
rect 4650 2148 4654 2204
rect 4654 2148 4710 2204
rect 4710 2148 4714 2204
rect 4650 2144 4714 2148
rect 4730 2204 4794 2208
rect 4730 2148 4734 2204
rect 4734 2148 4790 2204
rect 4790 2148 4794 2204
rect 4730 2144 4794 2148
rect 4810 2204 4874 2208
rect 4810 2148 4814 2204
rect 4814 2148 4870 2204
rect 4870 2148 4874 2204
rect 4810 2144 4874 2148
<< metal4 >>
rect 1848 7104 2168 7664
rect 1848 7040 1856 7104
rect 1920 7040 1936 7104
rect 2000 7040 2016 7104
rect 2080 7040 2096 7104
rect 2160 7040 2168 7104
rect 1848 6779 2168 7040
rect 1848 6543 1890 6779
rect 2126 6543 2168 6779
rect 1848 6016 2168 6543
rect 1848 5952 1856 6016
rect 1920 5952 1936 6016
rect 2000 5952 2016 6016
rect 2080 5952 2096 6016
rect 2160 5952 2168 6016
rect 1848 4966 2168 5952
rect 1848 4928 1890 4966
rect 2126 4928 2168 4966
rect 1848 4864 1856 4928
rect 2160 4864 2168 4928
rect 1848 4730 1890 4864
rect 2126 4730 2168 4864
rect 1848 3840 2168 4730
rect 1848 3776 1856 3840
rect 1920 3776 1936 3840
rect 2000 3776 2016 3840
rect 2080 3776 2096 3840
rect 2160 3776 2168 3840
rect 1848 3152 2168 3776
rect 1848 2916 1890 3152
rect 2126 2916 2168 3152
rect 1848 2752 2168 2916
rect 1848 2688 1856 2752
rect 1920 2688 1936 2752
rect 2000 2688 2016 2752
rect 2080 2688 2096 2752
rect 2160 2688 2168 2752
rect 1848 2128 2168 2688
rect 2753 7648 3074 7664
rect 2753 7584 2761 7648
rect 2825 7584 2841 7648
rect 2905 7584 2921 7648
rect 2985 7584 3001 7648
rect 3065 7584 3074 7648
rect 2753 6560 3074 7584
rect 2753 6496 2761 6560
rect 2825 6496 2841 6560
rect 2905 6496 2921 6560
rect 2985 6496 3001 6560
rect 3065 6496 3074 6560
rect 2753 5872 3074 6496
rect 2753 5636 2795 5872
rect 3031 5636 3074 5872
rect 2753 5472 3074 5636
rect 2753 5408 2761 5472
rect 2825 5408 2841 5472
rect 2905 5408 2921 5472
rect 2985 5408 3001 5472
rect 3065 5408 3074 5472
rect 2753 4384 3074 5408
rect 2753 4320 2761 4384
rect 2825 4320 2841 4384
rect 2905 4320 2921 4384
rect 2985 4320 3001 4384
rect 3065 4320 3074 4384
rect 2753 4059 3074 4320
rect 2753 3823 2795 4059
rect 3031 3823 3074 4059
rect 2753 3296 3074 3823
rect 2753 3232 2761 3296
rect 2825 3232 2841 3296
rect 2905 3232 2921 3296
rect 2985 3232 3001 3296
rect 3065 3232 3074 3296
rect 2753 2208 3074 3232
rect 2753 2144 2761 2208
rect 2825 2144 2841 2208
rect 2905 2144 2921 2208
rect 2985 2144 3001 2208
rect 3065 2144 3074 2208
rect 2753 2128 3074 2144
rect 3658 7104 3978 7664
rect 3658 7040 3666 7104
rect 3730 7040 3746 7104
rect 3810 7040 3826 7104
rect 3890 7040 3906 7104
rect 3970 7040 3978 7104
rect 3658 6779 3978 7040
rect 3658 6543 3700 6779
rect 3936 6543 3978 6779
rect 3658 6016 3978 6543
rect 3658 5952 3666 6016
rect 3730 5952 3746 6016
rect 3810 5952 3826 6016
rect 3890 5952 3906 6016
rect 3970 5952 3978 6016
rect 3658 4966 3978 5952
rect 3658 4928 3700 4966
rect 3936 4928 3978 4966
rect 3658 4864 3666 4928
rect 3970 4864 3978 4928
rect 3658 4730 3700 4864
rect 3936 4730 3978 4864
rect 3658 3840 3978 4730
rect 3658 3776 3666 3840
rect 3730 3776 3746 3840
rect 3810 3776 3826 3840
rect 3890 3776 3906 3840
rect 3970 3776 3978 3840
rect 3658 3152 3978 3776
rect 3658 2916 3700 3152
rect 3936 2916 3978 3152
rect 3658 2752 3978 2916
rect 3658 2688 3666 2752
rect 3730 2688 3746 2752
rect 3810 2688 3826 2752
rect 3890 2688 3906 2752
rect 3970 2688 3978 2752
rect 3658 2128 3978 2688
rect 4562 7648 4883 7664
rect 4562 7584 4570 7648
rect 4634 7584 4650 7648
rect 4714 7584 4730 7648
rect 4794 7584 4810 7648
rect 4874 7584 4883 7648
rect 4562 6560 4883 7584
rect 4562 6496 4570 6560
rect 4634 6496 4650 6560
rect 4714 6496 4730 6560
rect 4794 6496 4810 6560
rect 4874 6496 4883 6560
rect 4562 5872 4883 6496
rect 4562 5636 4604 5872
rect 4840 5636 4883 5872
rect 4562 5472 4883 5636
rect 4562 5408 4570 5472
rect 4634 5408 4650 5472
rect 4714 5408 4730 5472
rect 4794 5408 4810 5472
rect 4874 5408 4883 5472
rect 4562 4384 4883 5408
rect 4562 4320 4570 4384
rect 4634 4320 4650 4384
rect 4714 4320 4730 4384
rect 4794 4320 4810 4384
rect 4874 4320 4883 4384
rect 4562 4059 4883 4320
rect 4562 3823 4604 4059
rect 4840 3823 4883 4059
rect 4562 3296 4883 3823
rect 4562 3232 4570 3296
rect 4634 3232 4650 3296
rect 4714 3232 4730 3296
rect 4794 3232 4810 3296
rect 4874 3232 4883 3296
rect 4562 2208 4883 3232
rect 4562 2144 4570 2208
rect 4634 2144 4650 2208
rect 4714 2144 4730 2208
rect 4794 2144 4810 2208
rect 4874 2144 4883 2208
rect 4562 2128 4883 2144
rect 5467 7104 5787 7664
rect 5467 7040 5475 7104
rect 5539 7040 5555 7104
rect 5619 7040 5635 7104
rect 5699 7040 5715 7104
rect 5779 7040 5787 7104
rect 5467 6779 5787 7040
rect 5467 6543 5509 6779
rect 5745 6543 5787 6779
rect 5467 6016 5787 6543
rect 5467 5952 5475 6016
rect 5539 5952 5555 6016
rect 5619 5952 5635 6016
rect 5699 5952 5715 6016
rect 5779 5952 5787 6016
rect 5467 4966 5787 5952
rect 5467 4928 5509 4966
rect 5745 4928 5787 4966
rect 5467 4864 5475 4928
rect 5779 4864 5787 4928
rect 5467 4730 5509 4864
rect 5745 4730 5787 4864
rect 5467 3840 5787 4730
rect 5467 3776 5475 3840
rect 5539 3776 5555 3840
rect 5619 3776 5635 3840
rect 5699 3776 5715 3840
rect 5779 3776 5787 3840
rect 5467 3152 5787 3776
rect 5467 2916 5509 3152
rect 5745 2916 5787 3152
rect 5467 2752 5787 2916
rect 5467 2688 5475 2752
rect 5539 2688 5555 2752
rect 5619 2688 5635 2752
rect 5699 2688 5715 2752
rect 5779 2688 5787 2752
rect 5467 2128 5787 2688
<< via4 >>
rect 1890 6543 2126 6779
rect 1890 4928 2126 4966
rect 1890 4864 1920 4928
rect 1920 4864 1936 4928
rect 1936 4864 2000 4928
rect 2000 4864 2016 4928
rect 2016 4864 2080 4928
rect 2080 4864 2096 4928
rect 2096 4864 2126 4928
rect 1890 4730 2126 4864
rect 1890 2916 2126 3152
rect 2795 5636 3031 5872
rect 2795 3823 3031 4059
rect 3700 6543 3936 6779
rect 3700 4928 3936 4966
rect 3700 4864 3730 4928
rect 3730 4864 3746 4928
rect 3746 4864 3810 4928
rect 3810 4864 3826 4928
rect 3826 4864 3890 4928
rect 3890 4864 3906 4928
rect 3906 4864 3936 4928
rect 3700 4730 3936 4864
rect 3700 2916 3936 3152
rect 4604 5636 4840 5872
rect 4604 3823 4840 4059
rect 5509 6543 5745 6779
rect 5509 4928 5745 4966
rect 5509 4864 5539 4928
rect 5539 4864 5555 4928
rect 5555 4864 5619 4928
rect 5619 4864 5635 4928
rect 5635 4864 5699 4928
rect 5699 4864 5715 4928
rect 5715 4864 5745 4928
rect 5509 4730 5745 4864
rect 5509 2916 5745 3152
<< metal5 >>
rect 1104 6779 6532 6821
rect 1104 6543 1890 6779
rect 2126 6543 3700 6779
rect 3936 6543 5509 6779
rect 5745 6543 6532 6779
rect 1104 6501 6532 6543
rect 1104 5872 6532 5915
rect 1104 5636 2795 5872
rect 3031 5636 4604 5872
rect 4840 5636 6532 5872
rect 1104 5594 6532 5636
rect 1104 4966 6532 5008
rect 1104 4730 1890 4966
rect 2126 4730 3700 4966
rect 3936 4730 5509 4966
rect 5745 4730 6532 4966
rect 1104 4688 6532 4730
rect 1104 4059 6532 4101
rect 1104 3823 2795 4059
rect 3031 3823 4604 4059
rect 4840 3823 6532 4059
rect 1104 3781 6532 3823
rect 1104 3152 6532 3195
rect 1104 2916 1890 3152
rect 2126 2916 3700 3152
rect 3936 2916 5509 3152
rect 5745 2916 6532 3152
rect 1104 2874 6532 2916
use sky130_fd_sc_hd__decap_12  FILLER_0_3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1644511149
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_29
timestamp 1644511149
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_41
timestamp 1644511149
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1644511149
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1644511149
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1644511149
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1644511149
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1644511149
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1644511149
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1644511149
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1644511149
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_29
timestamp 1644511149
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_41
timestamp 1644511149
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_53
timestamp 1644511149
transform 1 0 5980 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1644511149
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1644511149
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1644511149
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1644511149
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1644511149
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1644511149
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1644511149
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1644511149
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1644511149
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_29
timestamp 1644511149
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_41
timestamp 1644511149
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_53
timestamp 1644511149
transform 1 0 5980 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1644511149
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1644511149
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1644511149
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_39 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 4692 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_47 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5428 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_52
timestamp 1644511149
transform 1 0 5888 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1644511149
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1644511149
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1644511149
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_29
timestamp 1644511149
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_41
timestamp 1644511149
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_53
timestamp 1644511149
transform 1 0 5980 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1644511149
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1644511149
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1644511149
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1644511149
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1644511149
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1644511149
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1644511149
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1644511149
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1644511149
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_29
timestamp 1644511149
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_41
timestamp 1644511149
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_53
timestamp 1644511149
transform 1 0 5980 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_6
timestamp 1644511149
transform 1 0 1656 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_18
timestamp 1644511149
transform 1 0 2760 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_26
timestamp 1644511149
transform 1 0 3496 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_29
timestamp 1644511149
transform 1 0 3772 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_41
timestamp 1644511149
transform 1 0 4876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_53
timestamp 1644511149
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1644511149
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1644511149
transform -1 0 6532 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1644511149
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1644511149
transform -1 0 6532 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1644511149
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1644511149
transform -1 0 6532 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1644511149
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1644511149
transform -1 0 6532 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1644511149
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1644511149
transform -1 0 6532 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1644511149
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1644511149
transform -1 0 6532 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1644511149
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1644511149
transform -1 0 6532 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1644511149
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1644511149
transform -1 0 6532 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1644511149
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1644511149
transform -1 0 6532 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1644511149
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1644511149
transform -1 0 6532 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_20 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_21
timestamp 1644511149
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_22
timestamp 1644511149
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_23
timestamp 1644511149
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_24
timestamp 1644511149
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_25
timestamp 1644511149
transform 1 0 3680 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _0__1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 1656 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1__2
timestamp 1644511149
transform 1 0 5612 0 -1 5440
box -38 -48 314 592
<< labels >>
rlabel metal5 s 1104 3781 6532 4101 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 5595 6532 5915 6 VGND
port 0 nsew ground input
rlabel metal4 s 2754 2128 3074 7664 6 VGND
port 0 nsew ground input
rlabel metal4 s 4563 2128 4883 7664 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 2875 6532 3195 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 4688 6532 5008 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 6501 6532 6821 6 VPWR
port 1 nsew power input
rlabel metal4 s 1848 2128 2168 7664 6 VPWR
port 1 nsew power input
rlabel metal4 s 3658 2128 3978 7664 6 VPWR
port 1 nsew power input
rlabel metal4 s 5467 2128 5787 7664 6 VPWR
port 1 nsew power input
rlabel metal3 s 0 2456 800 2576 6 avdd
port 2 nsew signal input
rlabel metal3 s 0 7352 800 7472 6 avss
port 3 nsew signal input
rlabel metal2 s 4802 9032 4858 9832 6 clk
port 4 nsew signal input
rlabel metal2 s 6734 0 6790 800 6 cvdd
port 5 nsew signal input
rlabel metal2 s 4802 0 4858 800 6 cvss
port 6 nsew signal input
rlabel metal2 s 2870 0 2926 800 6 dvdd
port 7 nsew signal input
rlabel metal2 s 938 0 994 800 6 dvss
port 8 nsew signal input
rlabel metal2 s 6734 9032 6790 9832 6 load
port 9 nsew signal input
rlabel metal2 s 938 9032 994 9832 6 out
port 10 nsew signal tristate
rlabel metal3 s 6888 8168 7688 8288 6 read
port 11 nsew signal input
rlabel metal2 s 2870 9032 2926 9832 6 ref
port 12 nsew signal input
rlabel metal3 s 6888 1640 7688 1760 6 s_in
port 13 nsew signal input
rlabel metal3 s 6888 4904 7688 5024 6 s_out
port 14 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 7688 9832
<< end >>
