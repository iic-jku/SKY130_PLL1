magic
tech sky130A
magscale 1 2
timestamp 1659939748
<< error_p >>
rect -461 151 -403 157
rect 403 151 461 157
rect -461 117 -449 151
rect 403 117 415 151
rect -461 111 -403 117
rect 403 111 461 117
<< nwell >>
rect -647 -289 647 289
<< pmos >>
rect -447 -70 -417 70
rect -351 -70 -321 70
rect -255 -70 -225 70
rect -159 -70 -129 70
rect -63 -70 -33 70
rect 33 -70 63 70
rect 129 -70 159 70
rect 225 -70 255 70
rect 321 -70 351 70
rect 417 -70 447 70
<< pdiff >>
rect -509 58 -447 70
rect -509 -58 -497 58
rect -463 -58 -447 58
rect -509 -70 -447 -58
rect -417 58 -351 70
rect -417 -58 -401 58
rect -367 -58 -351 58
rect -417 -70 -351 -58
rect -321 58 -255 70
rect -321 -58 -305 58
rect -271 -58 -255 58
rect -321 -70 -255 -58
rect -225 58 -159 70
rect -225 -58 -209 58
rect -175 -58 -159 58
rect -225 -70 -159 -58
rect -129 58 -63 70
rect -129 -58 -113 58
rect -79 -58 -63 58
rect -129 -70 -63 -58
rect -33 58 33 70
rect -33 -58 -17 58
rect 17 -58 33 58
rect -33 -70 33 -58
rect 63 58 129 70
rect 63 -58 79 58
rect 113 -58 129 58
rect 63 -70 129 -58
rect 159 58 225 70
rect 159 -58 175 58
rect 209 -58 225 58
rect 159 -70 225 -58
rect 255 58 321 70
rect 255 -58 271 58
rect 305 -58 321 58
rect 255 -70 321 -58
rect 351 58 417 70
rect 351 -58 367 58
rect 401 -58 417 58
rect 351 -70 417 -58
rect 447 58 509 70
rect 447 -58 463 58
rect 497 -58 509 58
rect 447 -70 509 -58
<< pdiffc >>
rect -497 -58 -463 58
rect -401 -58 -367 58
rect -305 -58 -271 58
rect -209 -58 -175 58
rect -113 -58 -79 58
rect -17 -58 17 58
rect 79 -58 113 58
rect 175 -58 209 58
rect 271 -58 305 58
rect 367 -58 401 58
rect 463 -58 497 58
<< nsubdiff >>
rect -611 219 -515 253
rect 515 219 611 253
rect -611 157 -577 219
rect 577 157 611 219
rect -611 -219 -577 -157
rect 577 -219 611 -157
rect -611 -253 -515 -219
rect 515 -253 611 -219
<< nsubdiffcont >>
rect -515 219 515 253
rect -611 -157 -577 157
rect 577 -157 611 157
rect -515 -253 515 -219
<< poly >>
rect -465 151 -399 167
rect -465 117 -449 151
rect -415 117 -399 151
rect -465 101 -399 117
rect 399 151 465 167
rect 399 117 415 151
rect 449 117 465 151
rect 399 101 465 117
rect -447 70 -417 101
rect -351 70 -321 96
rect -255 70 -225 96
rect -159 70 -129 96
rect -63 70 -33 96
rect 33 70 63 96
rect 129 70 159 96
rect 225 70 255 96
rect 321 70 351 96
rect 417 70 447 101
rect -447 -96 -417 -70
rect -351 -101 -321 -70
rect -255 -101 -225 -70
rect -159 -101 -129 -70
rect -63 -101 -33 -70
rect 33 -101 63 -70
rect 129 -101 159 -70
rect 225 -101 255 -70
rect 321 -101 351 -70
rect 417 -96 447 -70
rect -369 -117 369 -101
rect -369 -151 -353 -117
rect -319 -151 -257 -117
rect -223 -151 -161 -117
rect -127 -151 -65 -117
rect -31 -151 31 -117
rect 65 -151 127 -117
rect 161 -151 223 -117
rect 257 -151 319 -117
rect 353 -151 369 -117
rect -369 -167 369 -151
<< polycont >>
rect -449 117 -415 151
rect 415 117 449 151
rect -353 -151 -319 -117
rect -257 -151 -223 -117
rect -161 -151 -127 -117
rect -65 -151 -31 -117
rect 31 -151 65 -117
rect 127 -151 161 -117
rect 223 -151 257 -117
rect 319 -151 353 -117
<< locali >>
rect -611 219 -515 253
rect 515 219 611 253
rect -611 157 -577 219
rect 577 157 611 219
rect -465 117 -449 151
rect -415 117 -399 151
rect 399 117 415 151
rect 449 117 465 151
rect -497 58 -463 74
rect -497 -74 -463 -58
rect -401 58 -367 74
rect -401 -74 -367 -58
rect -305 58 -271 74
rect -305 -74 -271 -58
rect -209 58 -175 74
rect -209 -74 -175 -58
rect -113 58 -79 74
rect -113 -74 -79 -58
rect -17 58 17 74
rect -17 -74 17 -58
rect 79 58 113 74
rect 79 -74 113 -58
rect 175 58 209 74
rect 175 -74 209 -58
rect 271 58 305 74
rect 271 -74 305 -58
rect 367 58 401 74
rect 367 -74 401 -58
rect 463 58 497 74
rect 463 -74 497 -58
rect -369 -151 -353 -117
rect -319 -151 -257 -117
rect -223 -151 -161 -117
rect -127 -151 -65 -117
rect -31 -151 31 -117
rect 65 -151 127 -117
rect 161 -151 223 -117
rect 257 -151 319 -117
rect 353 -151 369 -117
rect -611 -219 -577 -157
rect 647 -58 717 12
rect 577 -219 611 -157
rect -611 -253 -515 -219
rect 515 -253 611 -219
<< viali >>
rect -449 117 -415 151
rect 415 117 449 151
rect -497 -58 -463 58
rect -401 -58 -367 58
rect -305 -58 -271 58
rect -209 -58 -175 58
rect -113 -58 -79 58
rect -17 -58 17 58
rect 79 -58 113 58
rect 175 -58 209 58
rect 271 -58 305 58
rect 367 -58 401 58
rect 463 -58 497 58
rect -353 -151 -319 -117
rect -257 -151 -223 -117
rect -161 -151 -127 -117
rect -65 -151 -31 -117
rect 31 -151 65 -117
rect 127 -151 161 -117
rect 223 -151 257 -117
rect 319 -151 353 -117
<< metal1 >>
rect -461 151 -403 157
rect -461 117 -449 151
rect -415 117 -403 151
rect -461 111 -403 117
rect 403 151 461 157
rect 403 117 415 151
rect 449 117 461 151
rect 403 111 461 117
rect -511 61 -449 70
rect -511 9 -506 61
rect -454 9 -449 61
rect -511 0 -497 9
rect -503 -58 -497 0
rect -463 0 -449 9
rect -415 61 -353 70
rect -415 9 -410 61
rect -358 9 -353 61
rect -415 0 -401 9
rect -463 -58 -457 0
rect -503 -70 -457 -58
rect -407 -58 -401 0
rect -367 0 -353 9
rect -311 58 -265 70
rect -311 0 -305 58
rect -367 -58 -361 0
rect -407 -70 -361 -58
rect -319 -9 -305 0
rect -271 0 -265 58
rect -223 61 -161 70
rect -223 9 -218 61
rect -166 9 -161 61
rect -223 0 -209 9
rect -271 -9 -257 0
rect -319 -61 -314 -9
rect -262 -61 -257 -9
rect -319 -70 -257 -61
rect -215 -58 -209 0
rect -175 0 -161 9
rect -119 58 -73 70
rect -119 0 -113 58
rect -175 -58 -169 0
rect -215 -70 -169 -58
rect -127 -9 -113 0
rect -79 0 -73 58
rect -31 61 31 70
rect -31 9 -26 61
rect 26 9 31 61
rect -31 0 -17 9
rect -79 -9 -65 0
rect -127 -61 -122 -9
rect -70 -61 -65 -9
rect -127 -70 -65 -61
rect -23 -58 -17 0
rect 17 0 31 9
rect 73 58 119 70
rect 73 0 79 58
rect 17 -58 23 0
rect -23 -70 23 -58
rect 65 -9 79 0
rect 113 0 119 58
rect 161 61 223 70
rect 161 9 166 61
rect 218 9 223 61
rect 161 0 175 9
rect 113 -9 127 0
rect 65 -61 70 -9
rect 122 -61 127 -9
rect 65 -70 127 -61
rect 169 -58 175 0
rect 209 0 223 9
rect 265 58 311 70
rect 265 0 271 58
rect 209 -58 215 0
rect 169 -70 215 -58
rect 257 -9 271 0
rect 305 0 311 58
rect 353 61 415 70
rect 353 9 358 61
rect 410 9 415 61
rect 353 0 367 9
rect 305 -9 319 0
rect 257 -61 262 -9
rect 314 -61 319 -9
rect 257 -70 319 -61
rect 361 -58 367 0
rect 401 0 415 9
rect 449 61 511 70
rect 449 9 454 61
rect 506 9 511 61
rect 449 0 463 9
rect 401 -58 407 0
rect 361 -70 407 -58
rect 457 -58 463 0
rect 497 0 511 9
rect 497 -58 503 0
rect 457 -70 503 -58
rect -365 -117 -307 -111
rect -269 -117 -211 -111
rect -173 -117 -115 -111
rect -77 -117 -19 -111
rect 19 -117 77 -111
rect 115 -117 173 -111
rect 211 -117 269 -111
rect 307 -117 365 -111
rect -365 -151 -353 -117
rect -319 -151 -257 -117
rect -223 -151 -161 -117
rect -127 -151 -65 -117
rect -31 -151 31 -117
rect 65 -151 127 -117
rect 161 -151 223 -117
rect 257 -151 319 -117
rect 353 -151 365 -117
rect -365 -157 -307 -151
rect -269 -157 -211 -151
rect -173 -157 -115 -151
rect -77 -157 -19 -151
rect 19 -157 77 -151
rect 115 -157 173 -151
rect 211 -157 269 -151
rect 307 -157 365 -151
<< via1 >>
rect -506 58 -454 61
rect -506 9 -497 58
rect -497 9 -463 58
rect -463 9 -454 58
rect -410 58 -358 61
rect -410 9 -401 58
rect -401 9 -367 58
rect -367 9 -358 58
rect -218 58 -166 61
rect -218 9 -209 58
rect -209 9 -175 58
rect -175 9 -166 58
rect -314 -58 -305 -9
rect -305 -58 -271 -9
rect -271 -58 -262 -9
rect -314 -61 -262 -58
rect -26 58 26 61
rect -26 9 -17 58
rect -17 9 17 58
rect 17 9 26 58
rect -122 -58 -113 -9
rect -113 -58 -79 -9
rect -79 -58 -70 -9
rect -122 -61 -70 -58
rect 166 58 218 61
rect 166 9 175 58
rect 175 9 209 58
rect 209 9 218 58
rect 70 -58 79 -9
rect 79 -58 113 -9
rect 113 -58 122 -9
rect 70 -61 122 -58
rect 358 58 410 61
rect 358 9 367 58
rect 367 9 401 58
rect 401 9 410 58
rect 262 -58 271 -9
rect 271 -58 305 -9
rect 305 -58 314 -9
rect 262 -61 314 -58
rect 454 58 506 61
rect 454 9 463 58
rect 463 9 497 58
rect 497 9 506 58
<< metal2 >>
rect -517 63 -347 72
rect -517 7 -508 63
rect -452 7 -412 63
rect -356 7 -347 63
rect -517 -2 -347 7
rect -229 63 -155 72
rect -229 7 -220 63
rect -164 7 -155 63
rect -319 -9 -257 0
rect -229 -2 -155 7
rect -37 63 37 72
rect -37 7 -28 63
rect 28 7 37 63
rect -319 -61 -314 -9
rect -262 -36 -257 -9
rect -127 -9 -65 0
rect -37 -2 37 7
rect 155 63 229 72
rect 155 7 164 63
rect 220 7 229 63
rect -127 -36 -122 -9
rect -262 -61 -122 -36
rect -70 -36 -65 -9
rect 65 -9 127 0
rect 155 -2 229 7
rect 347 63 517 72
rect 347 7 356 63
rect 412 7 452 63
rect 508 7 517 63
rect 65 -36 70 -9
rect -70 -61 70 -36
rect 122 -36 127 -9
rect 257 -9 319 0
rect 347 -2 517 7
rect 257 -36 262 -9
rect 122 -61 262 -36
rect 314 -61 319 -9
rect -319 -70 319 -61
<< via2 >>
rect -508 61 -452 63
rect -508 9 -506 61
rect -506 9 -454 61
rect -454 9 -452 61
rect -508 7 -452 9
rect -412 61 -356 63
rect -412 9 -410 61
rect -410 9 -358 61
rect -358 9 -356 61
rect -412 7 -356 9
rect -220 61 -164 63
rect -220 9 -218 61
rect -218 9 -166 61
rect -166 9 -164 61
rect -220 7 -164 9
rect -28 61 28 63
rect -28 9 -26 61
rect -26 9 26 61
rect 26 9 28 61
rect -28 7 28 9
rect 164 61 220 63
rect 164 9 166 61
rect 166 9 218 61
rect 218 9 220 61
rect 164 7 220 9
rect 356 61 412 63
rect 356 9 358 61
rect 358 9 410 61
rect 410 9 412 61
rect 356 7 412 9
rect 452 61 508 63
rect 452 9 454 61
rect 454 9 506 61
rect 506 9 508 61
rect 452 7 508 9
<< metal3 >>
rect -517 70 -347 72
rect -229 70 -155 72
rect -37 70 37 72
rect 155 70 229 72
rect 347 70 517 72
rect -517 63 517 70
rect -517 7 -508 63
rect -452 7 -412 63
rect -356 10 -220 63
rect -356 7 -347 10
rect -517 -2 -347 7
rect -229 7 -220 10
rect -164 10 -28 63
rect -164 7 -155 10
rect -229 -2 -155 7
rect -37 7 -28 10
rect 28 10 164 63
rect 28 7 37 10
rect -37 -2 37 7
rect 155 7 164 10
rect 220 10 356 63
rect 220 7 229 10
rect 155 -2 229 7
rect 347 7 356 10
rect 412 7 452 63
rect 508 7 517 63
rect 347 -2 517 7
<< properties >>
string FIXED_BBOX -594 -236 594 236
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.7 l 0.15 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
