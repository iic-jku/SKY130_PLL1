magic
tech sky130A
magscale 1 2
timestamp 1660928070
<< pwell >>
rect -359 -280 359 280
<< nmos >>
rect -159 -70 -129 70
rect -63 -70 -33 70
rect 33 -70 63 70
rect 129 -70 159 70
<< ndiff >>
rect -221 58 -159 70
rect -221 -58 -209 58
rect -175 -58 -159 58
rect -221 -70 -159 -58
rect -129 58 -63 70
rect -129 -58 -113 58
rect -79 -58 -63 58
rect -129 -70 -63 -58
rect -33 58 33 70
rect -33 -58 -17 58
rect 17 -58 33 58
rect -33 -70 33 -58
rect 63 58 129 70
rect 63 -58 79 58
rect 113 -58 129 58
rect 63 -70 129 -58
rect 159 58 221 70
rect 159 -58 175 58
rect 209 -58 221 58
rect 159 -70 221 -58
<< ndiffc >>
rect -209 -58 -175 58
rect -113 -58 -79 58
rect -17 -58 17 58
rect 79 -58 113 58
rect 175 -58 209 58
<< psubdiff >>
rect -323 210 -227 244
rect 227 210 323 244
rect -323 148 -289 210
rect 289 148 323 210
rect -323 -210 -289 -148
rect 289 -210 323 -148
rect -323 -244 -227 -210
rect 227 -244 323 -210
<< psubdiffcont >>
rect -227 210 227 244
rect -323 -148 -289 148
rect 289 -148 323 148
rect -227 -244 227 -210
<< poly >>
rect -177 142 -111 158
rect -177 108 -161 142
rect -127 108 -111 142
rect -177 92 -111 108
rect 111 142 177 158
rect 111 108 127 142
rect 161 108 177 142
rect -159 70 -129 92
rect -63 70 -33 96
rect 33 70 63 96
rect 111 92 177 108
rect 129 70 159 92
rect -159 -96 -129 -70
rect -63 -92 -33 -70
rect 33 -92 63 -70
rect -81 -108 81 -92
rect 129 -96 159 -70
rect -81 -142 -65 -108
rect -31 -142 31 -108
rect 65 -142 81 -108
rect -81 -158 81 -142
<< polycont >>
rect -161 108 -127 142
rect 127 108 161 142
rect -65 -142 -31 -108
rect 31 -142 65 -108
<< locali >>
rect -323 210 -227 244
rect 227 210 323 244
rect -323 148 -289 210
rect 289 148 323 210
rect -177 108 -161 142
rect -127 108 -111 142
rect 111 108 127 142
rect 161 108 177 142
rect -209 58 -175 74
rect -209 -74 -175 -58
rect -113 58 -79 74
rect -113 -74 -79 -58
rect -17 58 17 74
rect -17 -74 17 -58
rect 79 58 113 74
rect 79 -74 113 -58
rect 175 58 209 74
rect 175 -74 209 -58
rect -81 -142 -65 -108
rect -31 -142 31 -108
rect 65 -142 81 -108
rect -323 -210 -289 -148
rect 289 -210 323 -148
rect -323 -244 -227 -210
rect 227 -244 323 -210
<< viali >>
rect -161 108 -127 142
rect 127 108 161 142
rect -209 -58 -175 58
rect -113 -58 -79 58
rect -17 -58 17 58
rect 79 -58 113 58
rect 175 -58 209 58
rect -65 -142 -31 -108
rect 31 -142 65 -108
<< metal1 >>
rect -173 142 -115 148
rect 115 142 173 148
rect -173 108 -161 142
rect -127 108 127 142
rect 161 108 173 142
rect -173 102 -115 108
rect 115 102 173 108
rect -215 58 -169 70
rect -215 0 -209 58
rect -221 -9 -209 0
rect -175 0 -169 58
rect -119 58 -73 70
rect -119 0 -113 58
rect -175 -9 -113 0
rect -79 0 -73 58
rect -29 61 29 70
rect -29 9 -26 61
rect 26 9 29 61
rect -29 0 -17 9
rect -79 -9 -67 0
rect -221 -61 -218 -9
rect -166 -61 -122 -9
rect -70 -61 -67 -9
rect -221 -70 -67 -61
rect -23 -58 -17 0
rect 17 0 29 9
rect 73 58 119 70
rect 73 0 79 58
rect 17 -58 23 0
rect -23 -70 23 -58
rect 67 -9 79 0
rect 113 0 119 58
rect 169 58 215 70
rect 169 0 175 58
rect 113 -9 175 0
rect 209 0 215 58
rect 209 -9 221 0
rect 67 -61 70 -9
rect 122 -61 166 -9
rect 218 -61 221 -9
rect 67 -70 221 -61
rect -77 -108 77 -102
rect -77 -142 -65 -108
rect -31 -142 31 -108
rect 65 -142 77 -108
rect -77 -148 77 -142
<< via1 >>
rect -26 58 26 61
rect -26 9 -17 58
rect -17 9 17 58
rect 17 9 26 58
rect -218 -58 -209 -9
rect -209 -58 -175 -9
rect -175 -58 -166 -9
rect -218 -61 -166 -58
rect -122 -58 -113 -9
rect -113 -58 -79 -9
rect -79 -58 -70 -9
rect -122 -61 -70 -58
rect 70 -58 79 -9
rect 79 -58 113 -9
rect 113 -58 122 -9
rect 70 -61 122 -58
rect 166 -58 175 -9
rect 175 -58 209 -9
rect 209 -58 218 -9
rect 166 -61 218 -58
<< metal2 >>
rect -29 61 29 70
rect -29 9 -26 61
rect 26 9 29 61
rect -29 0 29 9
rect -221 -9 -67 0
rect -221 -61 -218 -9
rect -166 -61 -122 -9
rect -70 -28 -67 -9
rect 67 -9 221 0
rect 67 -28 70 -9
rect -70 -61 70 -28
rect 122 -61 166 -9
rect 218 -61 221 -9
rect -221 -70 221 -61
<< properties >>
string FIXED_BBOX -306 -227 306 227
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.7 l 0.150 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
