magic
tech sky130A
magscale 1 2
timestamp 1668291684
<< metal1 >>
rect -47040 14593 26131 14600
rect -47040 14590 1633 14593
rect -47040 13809 -23014 14590
rect -22962 13809 -21577 14590
rect -21525 13809 -14442 14590
rect -14390 13809 1633 14590
rect 1815 13809 8716 14593
rect 8898 13809 26131 14593
rect -47040 13800 26131 13809
rect -47526 13590 26131 13600
rect -47526 12809 -22375 13590
rect -22323 12809 -21456 13590
rect -21404 12809 -13803 13590
rect -13751 12809 26131 13590
rect -47526 12800 26131 12809
rect -22705 12630 -22699 12682
rect -22647 12630 -22641 12682
rect 1256 11675 1456 12800
rect 1626 12654 1826 12660
rect 1626 11675 1826 12454
rect 8705 12654 8905 12660
rect 8705 11824 8905 12454
rect 9075 11824 9275 12800
rect -14127 10469 -14075 10475
rect -14127 10411 -14075 10417
rect -14122 10334 -14080 10411
rect -22705 9308 -22699 9360
rect -22647 9308 -22641 9360
rect -2889 9308 -2883 9360
rect -2831 9308 -2825 9360
rect -22694 8856 -22652 9308
rect -2877 9271 -2837 9308
rect -21756 8915 -21750 8967
rect -21698 8962 -21692 8967
rect -21698 8920 -21353 8962
rect -21698 8915 -21692 8920
rect -19182 8742 -19176 8794
rect -19124 8742 -19118 8794
rect -16914 7601 -16908 7653
rect -16856 7601 -16850 7653
rect -11235 6832 -10664 6847
rect -11235 6767 -11220 6832
rect -13154 6725 -11220 6767
rect -22699 6598 -22647 6604
rect -22647 6551 -21311 6593
rect -22699 6540 -22647 6546
rect -18102 5460 -16168 5530
rect -16210 5335 -16168 5460
rect -13154 5403 -13112 6725
rect -11235 6654 -11220 6725
rect -10678 6654 -10664 6832
rect -11235 6641 -10664 6654
rect 12016 4118 12022 4170
rect 12074 4118 12080 4170
rect -16023 3103 -16017 3169
rect -15951 3103 -15294 3169
rect 895 1500 1095 3552
rect 9469 1500 9669 3552
rect -48429 1490 1300 1500
rect -48429 1489 -12990 1490
rect -48429 709 -18196 1489
rect -18144 709 -12990 1489
rect -12938 709 1300 1490
rect -48429 700 1300 709
rect 2100 700 2106 1500
rect 8494 700 8500 1500
rect 9300 700 26131 1500
rect -48290 493 1300 500
rect -48290 489 915 493
rect -48290 488 -21577 489
rect -48290 -287 -45447 488
rect -45039 -287 -21577 488
rect -48290 -291 -21577 -287
rect -21525 -291 -18558 489
rect -18506 -291 -12726 489
rect -12674 -291 915 489
rect 1097 -291 1300 493
rect -48290 -300 1300 -291
rect 2100 -300 2106 500
rect 8494 -300 8500 500
rect 9300 493 26131 500
rect 9300 -291 9461 493
rect 9643 488 26131 493
rect 9643 -287 25191 488
rect 25599 -287 26131 488
rect 9643 -291 26131 -287
rect 9300 -300 26131 -291
rect 12445 -393 12515 -387
rect 12445 -538 12515 -463
rect -18372 -573 -18252 -558
rect -18372 -1111 -18358 -573
rect -18266 -1111 -18252 -573
rect -18372 -1128 -18252 -1111
rect -1340 -573 -770 -558
rect -1340 -1111 -1096 -573
rect -1004 -1111 -770 -573
rect -1340 -1128 -770 -1111
rect 4771 -2504 5763 -2408
rect 2818 -3741 2870 -3735
rect 5626 -3741 5678 -3735
rect 2737 -3787 2818 -3747
rect 4851 -3747 4857 -3741
rect 4811 -3787 4857 -3747
rect 4851 -3793 4857 -3787
rect 4909 -3793 4915 -3741
rect 5678 -3787 5724 -3747
rect 7647 -3791 7653 -3739
rect 7705 -3745 7711 -3739
rect 7705 -3785 7798 -3745
rect 7705 -3791 7711 -3785
rect 2818 -3799 2870 -3793
rect 5626 -3799 5678 -3793
rect -44044 -11174 -43474 -10604
rect -42408 -11174 -41838 -10604
rect -40772 -11174 -40202 -10604
rect -39136 -11174 -38566 -10604
rect -37500 -11174 -36930 -10604
rect -35864 -11174 -35294 -10604
rect -34228 -11174 -33658 -10604
rect -32592 -11174 -32022 -10604
rect -30054 -11174 -29484 -10604
rect -28418 -11174 -27848 -10604
rect -26782 -11174 -26212 -10604
rect -25146 -11174 -24576 -10604
rect -23510 -11174 -22940 -10604
rect -21874 -11174 -21304 -10604
rect -20238 -11174 -19668 -10604
rect -18602 -11174 -18032 -10604
rect -16064 -11174 -15494 -10604
rect -14428 -11174 -13858 -10604
rect -12792 -11174 -12222 -10604
rect -11156 -11174 -10586 -10604
rect -9520 -11174 -8950 -10604
rect -7884 -11174 -7314 -10604
rect -6248 -11174 -5678 -10604
rect -4612 -11174 -4042 -10604
rect -2976 -11174 -2406 -10604
rect -1340 -11174 -770 -10604
rect 12172 -11154 12742 -10584
rect 13808 -11154 14378 -10584
rect 15444 -11140 16014 -10584
rect 15443 -11154 16014 -11140
rect 17080 -11154 17650 -10584
rect 18716 -11135 19286 -10584
rect 18715 -11154 19286 -11135
rect 20352 -11136 20922 -10584
rect 20351 -11154 20922 -11136
rect 21988 -11154 22558 -10584
rect 23624 -11154 24194 -10584
rect -44044 -57797 -43944 -11174
rect -42407 -57507 -42307 -11174
rect -40772 -57217 -40672 -11174
rect -39135 -56927 -39035 -11174
rect -37500 -56637 -37400 -11174
rect -35864 -56347 -35764 -11174
rect -34227 -56057 -34127 -11174
rect -32591 -55767 -32491 -11174
rect -30054 -11288 -29954 -11174
rect -30054 -11399 -29954 -11388
rect -28417 -11299 -28317 -11174
rect -28417 -11405 -28317 -11399
rect -26782 -11299 -26682 -11174
rect -26782 -11405 -26682 -11399
rect -25145 -11299 -25045 -11174
rect -25145 -11405 -25045 -11399
rect -23510 -11299 -23410 -11174
rect -23510 -11405 -23410 -11399
rect -21874 -11299 -21774 -11174
rect -21874 -11405 -21774 -11399
rect -20237 -11299 -20137 -11174
rect -20237 -11405 -20137 -11399
rect -18601 -11299 -18501 -11174
rect -18601 -11405 -18501 -11399
rect -16065 -11678 -15965 -11174
rect -26420 -11778 -15965 -11678
rect -26420 -13641 -26320 -11778
rect -14428 -11968 -14328 -11174
rect -23476 -12068 -14328 -11968
rect -23476 -13602 -23376 -12068
rect -12793 -12258 -12693 -11174
rect -23476 -13708 -23376 -13702
rect -20540 -12358 -12693 -12258
rect -20540 -13634 -20440 -12358
rect -11156 -12548 -11056 -11174
rect -20540 -13740 -20440 -13734
rect -17587 -12648 -11056 -12548
rect -17587 -13644 -17487 -12648
rect -9521 -12838 -9421 -11174
rect -26420 -13747 -26320 -13741
rect -17587 -13750 -17487 -13744
rect -14651 -12938 -9421 -12838
rect -14651 -13650 -14551 -12938
rect -7885 -13128 -7785 -11174
rect -14651 -13756 -14551 -13750
rect -11704 -13228 -7785 -13128
rect -11704 -13650 -11604 -13228
rect -8762 -13628 -8662 -13622
rect -6248 -13628 -6148 -11174
rect -8662 -13728 -6148 -13628
rect -5817 -13631 -5717 -13625
rect -4612 -13631 -4512 -11174
rect -2976 -13508 -2876 -11174
rect -2976 -13514 -2773 -13508
rect -2976 -13614 -2873 -13514
rect -1340 -13511 -1240 -11174
rect 74 -13511 174 -13505
rect -1340 -13611 74 -13511
rect -2873 -13620 -2773 -13614
rect 74 -13617 174 -13611
rect -8762 -13734 -8662 -13728
rect -5717 -13731 -4512 -13631
rect -5817 -13737 -5717 -13731
rect -11704 -13756 -11604 -13750
rect 12171 -26970 12271 -11154
rect 12171 -27079 12177 -26970
rect 12265 -27079 12271 -26970
rect 12171 -27093 12271 -27079
rect 13808 -30642 13908 -11154
rect 13808 -30751 13814 -30642
rect 13902 -30751 13908 -30642
rect 13808 -30765 13908 -30751
rect 15443 -34314 15543 -11154
rect 15443 -34423 15449 -34314
rect 15537 -34423 15543 -34314
rect 15443 -34437 15543 -34423
rect 17080 -37986 17180 -11154
rect 17080 -38095 17086 -37986
rect 17174 -38095 17180 -37986
rect 17080 -38109 17180 -38095
rect 18715 -41658 18815 -11154
rect 18715 -41767 18721 -41658
rect 18809 -41767 18815 -41658
rect 18715 -41780 18815 -41767
rect 20351 -45330 20451 -11154
rect 20351 -45439 20357 -45330
rect 20445 -45439 20451 -45330
rect 20351 -45453 20451 -45439
rect 21988 -49002 22088 -11154
rect 21988 -49111 21994 -49002
rect 22082 -49111 22088 -49002
rect 21988 -49125 22088 -49111
rect 23624 -52674 23724 -11154
rect 23624 -52783 23630 -52674
rect 23718 -52783 23724 -52674
rect 23624 -52797 23724 -52783
rect -26701 -55767 -26601 -55761
rect -32591 -55867 -26701 -55767
rect -26701 -55873 -26601 -55867
rect -23940 -56057 -23840 -56051
rect -34227 -56157 -23940 -56057
rect -23940 -56163 -23840 -56157
rect -21176 -56347 -21076 -56341
rect -35864 -56447 -21176 -56347
rect -21176 -56453 -21076 -56447
rect -18424 -56637 -18324 -56631
rect -37500 -56737 -18424 -56637
rect -18424 -56743 -18324 -56737
rect -15667 -56927 -15567 -56921
rect -39135 -57027 -15667 -56927
rect -15667 -57033 -15567 -57027
rect -12906 -57217 -12806 -57211
rect -40772 -57317 -12906 -57217
rect -12906 -57323 -12806 -57317
rect -10139 -57507 -10039 -57501
rect -42407 -57607 -10139 -57507
rect -10139 -57613 -10039 -57607
rect -7381 -57797 -7281 -57791
rect -44044 -57897 -7381 -57797
rect -7381 -57903 -7281 -57897
<< via1 >>
rect -23014 13809 -22962 14590
rect -21577 13809 -21525 14590
rect -14442 13809 -14390 14590
rect 1633 13809 1815 14593
rect 8716 13809 8898 14593
rect -22375 12809 -22323 13590
rect -21456 12809 -21404 13590
rect -13803 12809 -13751 13590
rect -22699 12630 -22647 12682
rect 1626 12454 1826 12654
rect 8705 12454 8905 12654
rect -14127 10417 -14075 10469
rect -22699 9308 -22647 9360
rect -2883 9308 -2831 9360
rect -21750 8915 -21698 8967
rect -19176 8742 -19124 8794
rect -16908 7601 -16856 7653
rect -22699 6546 -22647 6598
rect -11220 6654 -10678 6832
rect 12022 4118 12074 4170
rect -16017 3103 -15951 3169
rect -18196 709 -18144 1489
rect -12990 709 -12938 1490
rect 1300 700 2100 1500
rect 8500 700 9300 1500
rect -45447 -287 -45039 488
rect -21577 -291 -21525 489
rect -18558 -291 -18506 489
rect -12726 -291 -12674 489
rect 915 -291 1097 493
rect 1300 -300 2100 500
rect 8500 -300 9300 500
rect 9461 -291 9643 493
rect 25191 -287 25599 488
rect 12445 -463 12515 -393
rect -18358 -1111 -18266 -573
rect -1096 -1111 -1004 -573
rect 2818 -3793 2870 -3741
rect 4857 -3793 4909 -3741
rect 5626 -3793 5678 -3741
rect 7653 -3791 7705 -3739
rect -30054 -11388 -29954 -11288
rect -28417 -11399 -28317 -11299
rect -26782 -11399 -26682 -11299
rect -25145 -11399 -25045 -11299
rect -23510 -11399 -23410 -11299
rect -21874 -11399 -21774 -11299
rect -20237 -11399 -20137 -11299
rect -18601 -11399 -18501 -11299
rect -26420 -13741 -26320 -13641
rect -23476 -13702 -23376 -13602
rect -20540 -13734 -20440 -13634
rect -17587 -13744 -17487 -13644
rect -14651 -13750 -14551 -13650
rect -11704 -13750 -11604 -13650
rect -8762 -13728 -8662 -13628
rect -2873 -13614 -2773 -13514
rect 74 -13611 174 -13511
rect -5817 -13731 -5717 -13631
rect 12177 -27079 12265 -26970
rect 13814 -30751 13902 -30642
rect 15449 -34423 15537 -34314
rect 17086 -38095 17174 -37986
rect 18721 -41767 18809 -41658
rect 20357 -45439 20445 -45330
rect 21994 -49111 22082 -49002
rect 23630 -52783 23718 -52674
rect -26701 -55867 -26601 -55767
rect -23940 -56157 -23840 -56057
rect -21176 -56447 -21076 -56347
rect -18424 -56737 -18324 -56637
rect -15667 -57027 -15567 -56927
rect -12906 -57317 -12806 -57217
rect -10139 -57607 -10039 -57507
rect -7381 -57897 -7281 -57797
<< metal2 >>
rect -23023 14590 -22953 14600
rect -23023 13809 -23014 14590
rect -22962 13809 -22953 14590
rect -23023 12443 -22953 13809
rect -21586 14590 -21516 14600
rect -21586 13809 -21577 14590
rect -21525 13809 -21516 14590
rect -22384 13590 -22314 13600
rect -22384 12809 -22375 13590
rect -22323 12809 -22314 13590
rect -22699 12686 -22647 12688
rect -22712 12626 -22703 12686
rect -22643 12626 -22634 12686
rect -22699 12624 -22647 12626
rect -22384 12539 -22314 12809
rect -23023 8664 -22953 10802
rect -22694 10473 -22652 10515
rect -22712 10413 -22703 10473
rect -22643 10413 -22634 10473
rect -22699 9364 -22647 9366
rect -22712 9304 -22703 9364
rect -22643 9304 -22634 9364
rect -22699 9302 -22647 9304
rect -22384 8760 -22314 10610
rect -21750 8971 -21698 8973
rect -21763 8911 -21754 8971
rect -21694 8911 -21685 8971
rect -21750 8909 -21698 8911
rect -21586 7992 -21516 13809
rect -14451 14590 -14381 14600
rect -14451 13809 -14442 14590
rect -14390 13809 -14381 14590
rect -21465 13590 -21395 13600
rect -21465 12809 -21456 13590
rect -21404 12809 -21395 13590
rect -21465 8631 -21395 12809
rect -14451 10142 -14381 13809
rect 1626 14593 1826 14600
rect 1626 13809 1633 14593
rect 1815 13809 1826 14593
rect -13812 13590 -13742 13600
rect -13812 12809 -13803 13590
rect -13751 12809 -13742 13590
rect -14140 10413 -14131 10473
rect -14071 10413 -14062 10473
rect -13812 10238 -13742 12809
rect 1626 12654 1826 13809
rect 8705 14593 8905 14600
rect 8705 13809 8716 14593
rect 8898 13809 8905 14593
rect 8705 12654 8905 13809
rect 1620 12454 1626 12654
rect 1826 12454 1832 12654
rect 8699 12454 8705 12654
rect 8905 12454 8911 12654
rect -2883 9364 -2831 9366
rect -2896 9304 -2887 9364
rect -2827 9304 -2818 9364
rect -2883 9302 -2831 9304
rect -19176 8798 -19124 8800
rect -19189 8738 -19180 8798
rect -19120 8738 -19111 8798
rect -19176 8736 -19124 8738
rect 12146 8684 12155 8713
rect 12069 8642 12155 8684
rect 12146 8613 12155 8642
rect 12255 8613 12264 8713
rect -16908 7657 -16856 7659
rect -16921 7597 -16912 7657
rect -16852 7597 -16843 7657
rect -16908 7595 -16856 7597
rect -809 7090 -743 7156
rect -814 7085 -738 7090
rect -814 7019 -809 7085
rect -743 7019 -738 7085
rect -814 7014 -738 7019
rect -809 7010 -743 7014
rect -11235 6832 -10665 6849
rect -22694 6598 -22652 6736
rect -11235 6654 -11220 6832
rect -10678 6654 -10665 6832
rect -145 6800 -17 6809
rect -145 6690 -136 6800
rect -25 6775 -17 6800
rect -25 6715 -24 6775
rect -22 6715 -13 6775
rect -25 6690 -17 6715
rect -145 6681 -17 6690
rect -11235 6642 -10665 6654
rect 12146 6636 12155 6665
rect -22705 6546 -22699 6598
rect -22647 6546 -22641 6598
rect 12069 6594 12155 6636
rect 12146 6565 12155 6594
rect 12255 6565 12264 6665
rect -45460 488 -45028 500
rect -45460 -287 -45447 488
rect -45039 -287 -45028 488
rect -45460 -6464 -45028 -287
rect -21586 489 -21516 6292
rect 12146 4588 12155 4617
rect 12069 4546 12155 4588
rect 12146 4517 12155 4546
rect 12255 4517 12264 4617
rect 12022 4174 12074 4176
rect 12009 4114 12018 4174
rect 12078 4114 12087 4174
rect 12022 4112 12074 4114
rect -21586 -291 -21577 489
rect -21525 -291 -21516 489
rect -21586 -300 -21516 -291
rect -18567 3477 -16993 3547
rect -14141 3477 -12665 3547
rect -18567 489 -18497 3477
rect -16378 3298 -16369 3364
rect -16303 3298 -16088 3364
rect -16154 3169 -16088 3298
rect -16017 3169 -15951 3175
rect -16154 3103 -16017 3169
rect -16017 3097 -15951 3103
rect -18205 1489 -18135 2068
rect -18205 709 -18196 1489
rect -18144 709 -18135 1489
rect -18205 700 -18135 709
rect -12999 1490 -12929 2068
rect -12999 709 -12990 1490
rect -12938 709 -12929 1490
rect -12999 700 -12929 709
rect -18567 -291 -18558 489
rect -18506 -291 -18497 489
rect -18567 -300 -18497 -291
rect -12735 489 -12665 3477
rect -12735 -291 -12726 489
rect -12674 -291 -12665 489
rect -12735 -300 -12665 -291
rect 908 493 1108 3922
rect 1300 1500 2100 1506
rect 8500 1500 9300 1506
rect 1291 700 1300 1500
rect 2100 700 2109 1500
rect 8491 700 8500 1500
rect 9300 700 9309 1500
rect 1300 694 2100 700
rect 8500 694 9300 700
rect 1300 500 2100 506
rect 8500 500 9300 506
rect 908 -291 915 493
rect 1097 -291 1108 493
rect 908 -300 1108 -291
rect 1291 -300 1300 500
rect 2100 -300 2109 500
rect 8491 -300 8500 500
rect 9300 -300 9309 500
rect 9454 493 9654 3922
rect 9454 -291 9461 493
rect 9643 -291 9654 493
rect 9454 -300 9654 -291
rect 25178 488 25610 500
rect 25178 -287 25191 488
rect 25599 -287 25610 488
rect 1300 -306 2100 -300
rect 8500 -306 9300 -300
rect 12445 -393 12515 -384
rect 12439 -463 12445 -393
rect 12515 -463 12521 -393
rect 12445 -472 12515 -463
rect -18372 -573 -18252 -558
rect -18372 -1111 -18358 -573
rect -18266 -1111 -18252 -573
rect -18372 -1128 -18252 -1111
rect -1110 -573 -990 -558
rect -1110 -1111 -1096 -573
rect -1004 -1111 -990 -573
rect -1110 -1128 -990 -1111
rect 2814 -3737 2874 -3728
rect 4853 -3737 4913 -3728
rect 5622 -3737 5682 -3728
rect 7649 -3735 7709 -3726
rect 2812 -3793 2814 -3741
rect 2874 -3793 2876 -3741
rect 5620 -3793 5622 -3741
rect 5682 -3793 5684 -3741
rect 2814 -3806 2874 -3797
rect 4853 -3806 4913 -3797
rect 5622 -3806 5682 -3797
rect 7649 -3804 7709 -3795
rect 25178 -6444 25610 -287
rect -30060 -11388 -30054 -11288
rect -29954 -11388 -29948 -11288
rect -32018 -11488 -29954 -11388
rect -28423 -11399 -28417 -11299
rect -28317 -11399 -28311 -11299
rect -26788 -11399 -26782 -11299
rect -26682 -11399 -26676 -11299
rect -25151 -11399 -25145 -11299
rect -25045 -11399 -25039 -11299
rect -23516 -11399 -23510 -11299
rect -23410 -11399 -23404 -11299
rect -21880 -11399 -21874 -11299
rect -21774 -11399 -21768 -11299
rect -20243 -11399 -20237 -11299
rect -20137 -11399 -20131 -11299
rect -18607 -11399 -18601 -11299
rect -18501 -11399 -18495 -11299
rect -32018 -52673 -31918 -11488
rect -28417 -11678 -28317 -11399
rect -31728 -11778 -28317 -11678
rect -31728 -49001 -31628 -11778
rect -26782 -11968 -26682 -11399
rect -31438 -12068 -26682 -11968
rect -31438 -45329 -31338 -12068
rect -25145 -12258 -25045 -11399
rect -31148 -12358 -25045 -12258
rect -31148 -41657 -31048 -12358
rect -23510 -12548 -23410 -11399
rect -30858 -12648 -23410 -12548
rect -30858 -37985 -30758 -12648
rect -21874 -12838 -21774 -11399
rect -30568 -12938 -21774 -12838
rect -30568 -34313 -30468 -12938
rect -20237 -13128 -20137 -11399
rect -30278 -13228 -20137 -13128
rect -30278 -30641 -30178 -13228
rect -18601 -13418 -18501 -11399
rect -29988 -13518 -18501 -13418
rect -29988 -26969 -29888 -13518
rect -26426 -13741 -26420 -13641
rect -26320 -13741 -26314 -13641
rect -23482 -13702 -23476 -13602
rect -23376 -13702 -23370 -13602
rect -2879 -13614 -2873 -13514
rect -2773 -13614 -2767 -13514
rect 68 -13611 74 -13511
rect 174 -13611 180 -13511
rect -26402 -13889 -26346 -13741
rect -23458 -13863 -23402 -13702
rect -20546 -13734 -20540 -13634
rect -20440 -13734 -20434 -13634
rect -20514 -13889 -20458 -13734
rect -17593 -13744 -17587 -13644
rect -17487 -13744 -17481 -13644
rect -17570 -13863 -17514 -13744
rect -14657 -13750 -14651 -13650
rect -14551 -13750 -14545 -13650
rect -11710 -13750 -11704 -13650
rect -11604 -13750 -11598 -13650
rect -8768 -13728 -8762 -13628
rect -8662 -13728 -8656 -13628
rect -14626 -13863 -14570 -13750
rect -11682 -13863 -11626 -13750
rect -8738 -13871 -8682 -13728
rect -5823 -13731 -5817 -13631
rect -5717 -13731 -5711 -13631
rect -5794 -13863 -5738 -13731
rect -2850 -13863 -2794 -13614
rect 94 -13863 150 -13611
rect 3038 -13871 3094 -13536
rect 5982 -13863 6038 -13548
rect 8900 -13600 26051 -13500
rect 8926 -13863 8982 -13600
rect 12171 -26964 12271 -26955
rect -29988 -27079 -29984 -26969
rect -29892 -27079 -29888 -26969
rect -29988 -27094 -29888 -27079
rect 12162 -26970 12279 -26964
rect 12162 -27079 12177 -26970
rect 12265 -27079 12279 -26970
rect 12162 -27084 12279 -27079
rect 12171 -27093 12271 -27084
rect 13808 -30636 13908 -30627
rect -30278 -30751 -30274 -30641
rect -30182 -30751 -30178 -30641
rect -30278 -30766 -30178 -30751
rect 13799 -30642 13916 -30636
rect 13799 -30751 13814 -30642
rect 13902 -30751 13916 -30642
rect 13799 -30756 13916 -30751
rect 13808 -30765 13908 -30756
rect 15443 -34308 15543 -34299
rect -30568 -34423 -30564 -34313
rect -30472 -34423 -30468 -34313
rect -30568 -34438 -30468 -34423
rect 15434 -34314 15551 -34308
rect 15434 -34423 15449 -34314
rect 15537 -34423 15551 -34314
rect 15434 -34428 15551 -34423
rect 15443 -34437 15543 -34428
rect 17080 -37980 17180 -37971
rect -30858 -38095 -30854 -37985
rect -30762 -38095 -30758 -37985
rect -30858 -38110 -30758 -38095
rect 17071 -37986 17188 -37980
rect 17071 -38095 17086 -37986
rect 17174 -38095 17188 -37986
rect 17071 -38100 17188 -38095
rect 17080 -38109 17180 -38100
rect 18715 -41652 18815 -41643
rect -31148 -41767 -31144 -41657
rect -31052 -41767 -31048 -41657
rect -31148 -41782 -31048 -41767
rect 18706 -41658 18823 -41652
rect 18706 -41767 18721 -41658
rect 18809 -41767 18823 -41658
rect 18706 -41772 18823 -41767
rect 18715 -41781 18815 -41772
rect 20351 -45324 20451 -45315
rect -31438 -45439 -31434 -45329
rect -31342 -45439 -31338 -45329
rect -31438 -45454 -31338 -45439
rect 20342 -45330 20459 -45324
rect 20342 -45439 20357 -45330
rect 20445 -45439 20459 -45330
rect 20342 -45444 20459 -45439
rect 20351 -45453 20451 -45444
rect 21988 -48996 22088 -48987
rect -31728 -49111 -31724 -49001
rect -31632 -49111 -31628 -49001
rect -31728 -49126 -31628 -49111
rect 21979 -49002 22096 -48996
rect 21979 -49111 21994 -49002
rect 22082 -49111 22096 -49002
rect 21979 -49116 22096 -49111
rect 21988 -49125 22088 -49116
rect 23624 -52668 23724 -52659
rect -32018 -52783 -32014 -52673
rect -31922 -52783 -31918 -52673
rect -32018 -52798 -31918 -52783
rect 23615 -52674 23732 -52668
rect 23615 -52783 23630 -52674
rect 23718 -52783 23732 -52674
rect 23615 -52788 23732 -52783
rect 23624 -52797 23724 -52788
rect -26678 -54901 -26622 -54616
rect -23918 -54901 -23862 -54628
rect -21158 -54898 -21102 -54640
rect -18398 -54895 -18342 -54640
rect -26701 -55767 -26601 -54901
rect -26707 -55867 -26701 -55767
rect -26601 -55867 -26595 -55767
rect -23940 -56057 -23840 -54901
rect -23946 -56157 -23940 -56057
rect -23840 -56157 -23834 -56057
rect -21176 -56347 -21076 -54898
rect -21182 -56447 -21176 -56347
rect -21076 -56447 -21070 -56347
rect -18424 -56637 -18324 -54895
rect -15638 -54898 -15582 -54628
rect -12878 -54898 -12822 -54593
rect -18430 -56737 -18424 -56637
rect -18324 -56737 -18318 -56637
rect -15667 -56927 -15567 -54898
rect -15673 -57027 -15667 -56927
rect -15567 -57027 -15561 -56927
rect -12906 -57217 -12806 -54898
rect -10118 -54901 -10062 -54616
rect -7358 -54898 -7302 -54605
rect -4598 -54892 -4542 -54605
rect -1838 -54891 -1782 -54628
rect 922 -54890 978 -54628
rect -12912 -57317 -12906 -57217
rect -12806 -57317 -12800 -57217
rect -10139 -57507 -10039 -54901
rect -10145 -57607 -10139 -57507
rect -10039 -57607 -10033 -57507
rect -7381 -57797 -7281 -54898
rect -4622 -54901 -4522 -54892
rect -4622 -55010 -4522 -55001
rect -1860 -54900 -1760 -54891
rect -1860 -55009 -1760 -55000
rect 899 -54899 999 -54890
rect 3682 -54891 3738 -54628
rect 6442 -54891 6498 -54628
rect 9202 -54891 9258 -54628
rect 899 -55008 999 -54999
rect 3659 -54900 3759 -54891
rect 3659 -55009 3759 -55000
rect 6419 -54900 6519 -54891
rect 6419 -55009 6519 -55000
rect 9179 -54900 9279 -54891
rect 9179 -55009 9279 -55000
rect -7387 -57897 -7381 -57797
rect -7281 -57897 -7275 -57797
<< via2 >>
rect -22703 12682 -22643 12686
rect -22703 12630 -22699 12682
rect -22699 12630 -22647 12682
rect -22647 12630 -22643 12682
rect -22703 12626 -22643 12630
rect -22703 10413 -22643 10473
rect -22703 9360 -22643 9364
rect -22703 9308 -22699 9360
rect -22699 9308 -22647 9360
rect -22647 9308 -22643 9360
rect -22703 9304 -22643 9308
rect -21754 8967 -21694 8971
rect -21754 8915 -21750 8967
rect -21750 8915 -21698 8967
rect -21698 8915 -21694 8967
rect -21754 8911 -21694 8915
rect -14131 10469 -14071 10473
rect -14131 10417 -14127 10469
rect -14127 10417 -14075 10469
rect -14075 10417 -14071 10469
rect -14131 10413 -14071 10417
rect -2887 9360 -2827 9364
rect -2887 9308 -2883 9360
rect -2883 9308 -2831 9360
rect -2831 9308 -2827 9360
rect -2887 9304 -2827 9308
rect -19180 8794 -19120 8798
rect -19180 8742 -19176 8794
rect -19176 8742 -19124 8794
rect -19124 8742 -19120 8794
rect -19180 8738 -19120 8742
rect 12155 8613 12255 8713
rect -16912 7653 -16852 7657
rect -16912 7601 -16908 7653
rect -16908 7601 -16856 7653
rect -16856 7601 -16852 7653
rect -16912 7597 -16852 7601
rect -809 7019 -743 7085
rect -136 6690 -25 6800
rect 12155 6565 12255 6665
rect 12155 4517 12255 4617
rect 12018 4170 12078 4174
rect 12018 4118 12022 4170
rect 12022 4118 12074 4170
rect 12074 4118 12078 4170
rect 12018 4114 12078 4118
rect -16369 3298 -16303 3364
rect 1300 700 2100 1500
rect 8500 700 9300 1500
rect 1300 -300 2100 500
rect 8500 -300 9300 500
rect 12445 -463 12515 -393
rect -18358 -1111 -18266 -573
rect -1096 -1111 -1004 -573
rect 2814 -3741 2874 -3737
rect 4853 -3741 4913 -3737
rect 5622 -3741 5682 -3737
rect 7649 -3739 7709 -3735
rect 2814 -3793 2818 -3741
rect 2818 -3793 2870 -3741
rect 2870 -3793 2874 -3741
rect 4853 -3793 4857 -3741
rect 4857 -3793 4909 -3741
rect 4909 -3793 4913 -3741
rect 5622 -3793 5626 -3741
rect 5626 -3793 5678 -3741
rect 5678 -3793 5682 -3741
rect 7649 -3791 7653 -3739
rect 7653 -3791 7705 -3739
rect 7705 -3791 7709 -3739
rect 2814 -3797 2874 -3793
rect 4853 -3797 4913 -3793
rect 5622 -3797 5682 -3793
rect 7649 -3795 7709 -3791
rect -29984 -27079 -29892 -26969
rect 12177 -27079 12265 -26970
rect -30274 -30751 -30182 -30641
rect 13814 -30751 13902 -30642
rect -30564 -34423 -30472 -34313
rect 15449 -34423 15537 -34314
rect -30854 -38095 -30762 -37985
rect 17086 -38095 17174 -37986
rect -31144 -41767 -31052 -41657
rect 18721 -41767 18809 -41658
rect -31434 -45439 -31342 -45329
rect 20357 -45439 20445 -45330
rect -31724 -49111 -31632 -49001
rect 21994 -49111 22082 -49002
rect -32014 -52783 -31922 -52673
rect 23630 -52783 23718 -52674
rect -4622 -55001 -4522 -54901
rect -1860 -55000 -1760 -54900
rect 899 -54999 999 -54899
rect 3659 -55000 3759 -54900
rect 6419 -55000 6519 -54900
rect 9179 -55000 9279 -54900
<< metal3 >>
rect -22708 12686 -22638 12691
rect -24440 12626 -22703 12686
rect -22643 12626 -22638 12686
rect -22708 12621 -22638 12626
rect -22708 10473 -22638 10478
rect -14136 10473 -14066 10478
rect -22708 10413 -22703 10473
rect -22643 10413 -14131 10473
rect -14071 10413 -14066 10473
rect -22708 10408 -22638 10413
rect -14136 10408 -14066 10413
rect -22708 9366 -22638 9369
rect -2892 9366 -2822 9369
rect -22711 9302 -22705 9366
rect -22641 9364 -22635 9366
rect -2895 9364 -2889 9366
rect -22641 9304 -22551 9364
rect -2977 9304 -2889 9364
rect -22641 9302 -22635 9304
rect -2895 9302 -2889 9304
rect -2825 9302 -2819 9366
rect -22708 9299 -22638 9302
rect -2892 9299 -2822 9302
rect -21759 8971 -21689 8976
rect -21991 8911 -21754 8971
rect -21694 8911 -21689 8971
rect -21991 3376 -21931 8911
rect -21759 8906 -21689 8911
rect -19185 8798 -19115 8803
rect -29397 3276 -21931 3376
rect -21850 8738 -19180 8798
rect -19120 8738 -19115 8798
rect -29397 -23292 -29297 3276
rect -21850 2976 -21790 8738
rect -19185 8733 -19115 8738
rect 12150 8713 12260 8718
rect 12150 8613 12155 8713
rect 12255 8613 13715 8713
rect 12150 8608 12260 8613
rect -16917 7657 -16847 7662
rect -28997 2876 -21790 2976
rect -21709 7597 -16912 7657
rect -16852 7597 -16847 7657
rect -28997 -19620 -28897 2876
rect -21709 2576 -21649 7597
rect -16917 7592 -16847 7597
rect -814 7085 -738 7090
rect -814 7019 -809 7085
rect -743 7082 -738 7085
rect -743 7022 548 7082
rect -743 7019 -738 7022
rect -814 7014 -738 7019
rect -8027 6800 -17 6809
rect -8027 6690 -136 6800
rect -25 6690 -17 6800
rect -8027 6681 -17 6690
rect -16374 3364 -16298 3369
rect -28597 2476 -21649 2576
rect -18343 3298 -16369 3364
rect -16303 3298 -16298 3364
rect -28597 -15948 -28497 2476
rect -18343 -558 -18277 3298
rect -16374 3293 -16298 3298
rect -1081 -558 -1015 6681
rect 12150 6665 12260 6670
rect 12150 6565 12155 6665
rect 12255 6565 13315 6665
rect 12150 6560 12260 6565
rect 12150 4617 12260 4622
rect 12150 4517 12155 4617
rect 12255 4517 12915 4617
rect 12150 4512 12260 4517
rect 12013 4174 12515 4179
rect 12013 4114 12018 4174
rect 12078 4114 12515 4174
rect 12013 4109 12515 4114
rect 1295 1500 2105 1505
rect 8495 1500 9305 1505
rect 1295 700 1300 1500
rect 2100 700 8500 1500
rect 9300 700 9305 1500
rect 1295 695 2105 700
rect 8495 695 9305 700
rect 1295 500 2105 505
rect 8495 500 9305 505
rect 1295 -300 1300 500
rect 2100 -300 8500 500
rect 9300 -300 9305 500
rect 1295 -305 2105 -300
rect 8495 -305 9305 -300
rect 12445 -388 12515 4109
rect 12440 -393 12520 -388
rect 12440 -463 12445 -393
rect 12515 -463 12520 -393
rect 12440 -468 12520 -463
rect -18372 -573 -18252 -558
rect -18372 -1111 -18358 -573
rect -18266 -1111 -18252 -573
rect -18372 -1128 -18252 -1111
rect -1110 -573 -990 -558
rect -1110 -1111 -1096 -573
rect -1004 -1111 -990 -573
rect -1110 -1128 -990 -1111
rect 2809 -3737 2879 -3732
rect 2809 -3797 2814 -3737
rect 2874 -3797 2879 -3737
rect 2809 -3802 2879 -3797
rect 4848 -3737 4918 -3732
rect 4848 -3797 4853 -3737
rect 4913 -3797 4918 -3737
rect 4848 -3802 4918 -3797
rect 5617 -3737 5687 -3732
rect 5617 -3797 5622 -3737
rect 5682 -3797 5687 -3737
rect 5617 -3802 5687 -3797
rect 7644 -3735 7714 -3730
rect 7644 -3795 7649 -3735
rect 7709 -3795 7714 -3735
rect 7644 -3800 7714 -3795
rect 2814 -8680 2874 -3802
rect 4853 -8680 4913 -3802
rect 5622 -8680 5682 -3802
rect 7649 -8680 7709 -3800
rect 12815 -15948 12915 4517
rect -28597 -16068 -27956 -15948
rect 10553 -16068 12915 -15948
rect 13215 -19620 13315 6565
rect -28997 -19740 -27956 -19620
rect 10553 -19740 13315 -19620
rect 13615 -23292 13715 8613
rect -29397 -23412 -27956 -23292
rect 10506 -23412 13715 -23292
rect -29998 -26969 -27956 -26964
rect -29998 -27079 -29984 -26969
rect -29892 -27079 -27956 -26969
rect -29998 -27084 -27956 -27079
rect 10553 -26970 12286 -26964
rect 10553 -27079 12177 -26970
rect 12265 -27079 12286 -26970
rect 10553 -27084 12286 -27079
rect -30288 -30641 -27949 -30636
rect -30288 -30751 -30274 -30641
rect -30182 -30751 -27949 -30641
rect -30288 -30756 -27949 -30751
rect 10506 -30642 13923 -30636
rect 10506 -30751 13814 -30642
rect 13902 -30751 13923 -30642
rect 10506 -30756 13923 -30751
rect -30578 -34313 -27956 -34308
rect -30578 -34423 -30564 -34313
rect -30472 -34423 -27956 -34313
rect -30578 -34428 -27956 -34423
rect 10529 -34314 15558 -34308
rect 10529 -34423 15449 -34314
rect 15537 -34423 15558 -34314
rect 10529 -34428 15558 -34423
rect -30868 -37985 -27914 -37980
rect -30868 -38095 -30854 -37985
rect -30762 -38095 -27914 -37985
rect -30868 -38100 -27914 -38095
rect 10529 -37986 17195 -37980
rect 10529 -38095 17086 -37986
rect 17174 -38095 17195 -37986
rect 10529 -38100 17195 -38095
rect -31158 -41657 -27949 -41652
rect -31158 -41767 -31144 -41657
rect -31052 -41767 -27949 -41657
rect -31158 -41772 -27949 -41767
rect 10518 -41658 18830 -41652
rect 10518 -41767 18721 -41658
rect 18809 -41767 18830 -41658
rect 10518 -41772 18830 -41767
rect -31448 -45329 -27956 -45324
rect -31448 -45439 -31434 -45329
rect -31342 -45439 -27956 -45329
rect -31448 -45444 -27956 -45439
rect 10506 -45330 20466 -45324
rect 10506 -45439 20357 -45330
rect 20445 -45439 20466 -45330
rect 10506 -45444 20466 -45439
rect -31738 -49001 -27956 -48996
rect -31738 -49111 -31724 -49001
rect -31632 -49111 -27956 -49001
rect -31738 -49116 -27956 -49111
rect 10553 -49002 22103 -48996
rect 10553 -49111 21994 -49002
rect 22082 -49111 22103 -49002
rect 10553 -49116 22103 -49111
rect -32028 -52673 -27956 -52668
rect -32028 -52783 -32014 -52673
rect -31922 -52783 -27956 -52673
rect -32028 -52788 -27956 -52783
rect 10506 -52674 23739 -52668
rect 10506 -52783 23630 -52674
rect 23718 -52783 23739 -52674
rect 10506 -52788 23739 -52783
rect -4627 -54901 -4517 -54896
rect -4627 -55001 -4622 -54901
rect -4522 -55001 -4517 -54901
rect -4627 -55006 -4517 -55001
rect -1865 -54900 -1755 -54895
rect -1865 -55000 -1860 -54900
rect -1760 -55000 -1755 -54900
rect -1865 -55005 -1755 -55000
rect 894 -54899 1004 -54894
rect 894 -54999 899 -54899
rect 999 -54999 1004 -54899
rect 894 -55004 1004 -54999
rect 3654 -54900 3764 -54895
rect 3654 -55000 3659 -54900
rect 3759 -55000 3764 -54900
rect -4622 -58300 -4522 -55006
rect -1860 -58300 -1760 -55005
rect 899 -58300 999 -55004
rect 3654 -55005 3764 -55000
rect 6414 -54900 6524 -54895
rect 6414 -55000 6419 -54900
rect 6519 -55000 6524 -54900
rect 6414 -55005 6524 -55000
rect 9174 -54900 9284 -54895
rect 9174 -55000 9179 -54900
rect 9279 -55000 9284 -54900
rect 9174 -55005 9284 -55000
rect 3659 -58300 3759 -55005
rect 6419 -58300 6519 -55005
rect 9179 -58300 9279 -55005
<< via3 >>
rect -22705 9364 -22641 9366
rect -2889 9364 -2825 9366
rect -22705 9304 -22703 9364
rect -22703 9304 -22643 9364
rect -22643 9304 -22641 9364
rect -2889 9304 -2887 9364
rect -2887 9304 -2827 9364
rect -2827 9304 -2825 9364
rect -22705 9302 -22641 9304
rect -2889 9302 -2825 9304
<< metal4 >>
rect -22706 9366 -22640 9367
rect -22706 9364 -22705 9366
rect -22714 9304 -22705 9364
rect -22706 9302 -22705 9304
rect -22641 9364 -22640 9366
rect -2890 9366 -2824 9367
rect -2890 9364 -2889 9366
rect -22641 9304 -2889 9364
rect -22641 9302 -22640 9304
rect -22706 9301 -22640 9302
rect -2890 9302 -2889 9304
rect -2825 9302 -2824 9366
rect -2890 9301 -2824 9302
use d_ff_15  d_ff_15_0
timestamp 1668240031
transform 0 1 -1002 1 0 7173
box -98 -2224 2138 697
use full_vco_1  full_vco_1_0
timestamp 1668250571
transform 1 0 1247 0 1 3352
box -1329 -7488 10864 8523
use inv_buffer2  inv_buffer2_0
timestamp 1668240031
transform 0 1 2989 -1 0 -8970
box 0 0 2204 1138
use inv_buffer2  inv_buffer2_1
timestamp 1668240031
transform 0 -1 5265 -1 0 -8970
box 0 0 2204 1138
use inv_buffer2  inv_buffer2_2
timestamp 1668240031
transform 0 1 5265 -1 0 -8970
box 0 0 2204 1138
use inv_buffer2  inv_buffer2_3
timestamp 1668240031
transform 0 -1 7541 -1 0 -8970
box 0 0 2204 1138
use inv_buffer2  inv_buffer2_8
timestamp 1668240031
transform 0 1 -23233 -1 0 8898
box 0 0 2204 1138
use inv_buffer2  inv_buffer2_9
timestamp 1668240031
transform 0 1 -23193 -1 0 12677
box 0 0 2204 1138
use r2r_8  r2r_8_0
timestamp 1668290053
transform -1 0 25125 0 1 -10561
box -485 -593 13937 10023
use r2r_8  r2r_8_1
timestamp 1668290053
transform 1 0 -30985 0 1 -10581
box -485 -593 13937 10023
use r2r_8  r2r_8_2
timestamp 1668290053
transform 1 0 -44975 0 1 -10581
box -485 -593 13937 10023
use r2r_10  r2r_10_0
timestamp 1668290266
transform 1 0 -16995 0 1 -10581
box -485 -593 17209 10023
use slopebuf  slopebuf_0
timestamp 1668240031
transform 1 0 -21311 0 1 6012
box -866 -1740 4686 2950
use sspd  sspd_0
timestamp 1668291684
transform 0 1 -18419 -1 0 9251
box -1125 214 7472 5865
use voltage_control  voltage_control_0
timestamp 1668291684
transform 1 0 -82459 0 1 -4512
box 41052 6053 104762 89673
use wrapper  wrapper_0 wrapper/runs/RUN_2022.11.11_11.09.27/results/final/mag
timestamp 1668240031
transform 1 0 -28076 0 1 -54700
box 0 0 38749 40893
<< labels >>
rlabel metal1 -1340 -1128 -770 -558 0 vout
<< end >>
