magic
tech sky130A
magscale 1 2
timestamp 1668357910
<< metal1 >>
rect 1540 1436 1582 1528
rect 1801 1182 1871 1188
rect 1801 871 1871 1112
rect 1801 795 1871 801
rect 2440 1187 2510 1193
rect 2440 871 2510 1117
rect 2440 795 2510 801
rect 1540 -608 1582 -516
rect 1801 -864 1871 -858
rect 1801 -1164 1871 -934
rect 2440 -873 2510 -867
rect 2440 -1145 2510 -943
rect 2440 -1221 2510 -1215
rect 1801 -1240 1871 -1234
rect 1540 -2564 1582 -2522
<< via1 >>
rect 1801 1112 1871 1182
rect 1801 801 1871 871
rect 2440 1117 2510 1187
rect 2440 801 2510 871
rect 1801 -934 1871 -864
rect 1801 -1234 1871 -1164
rect 2440 -943 2510 -873
rect 2440 -1215 2510 -1145
<< metal2 >>
rect 1498 3019 1540 3061
rect 2720 3019 2762 3061
rect 1801 1182 1871 1708
rect 2440 1187 2510 1804
rect 1795 1112 1801 1182
rect 1871 1112 1877 1182
rect 2434 1117 2440 1187
rect 2510 1117 2516 1187
rect 1498 973 1540 1015
rect 2720 973 2762 1015
rect 1795 801 1801 871
rect 1871 801 1877 871
rect 2434 801 2440 871
rect 2510 801 2516 871
rect 1801 294 1871 801
rect 2440 197 2510 801
rect 1801 -864 1871 -336
rect 1795 -934 1801 -864
rect 1871 -934 1877 -864
rect 2440 -873 2510 -240
rect 2434 -943 2440 -873
rect 2510 -943 2516 -873
rect 1498 -1073 1540 -1031
rect 2720 -1073 2762 -1031
rect 1795 -1234 1801 -1164
rect 1871 -1234 1877 -1164
rect 2434 -1215 2440 -1145
rect 2510 -1215 2516 -1145
rect 1801 -1754 1871 -1234
rect 2440 -1850 2510 -1215
rect 2440 -2358 2510 -2288
rect 1801 -2455 1871 -2385
use tgate_1  tgate_1_0
timestamp 1668357910
transform 1 0 1801 0 1 2480
box -261 -952 919 1138
use tgate_1  tgate_1_1
timestamp 1668357910
transform 1 0 1801 0 1 434
box -261 -952 919 1138
use tgate_1  tgate_1_2
timestamp 1668357910
transform 1 0 1801 0 1 -1612
box -261 -952 919 1138
<< labels >>
rlabel metal2 2720 3019 2762 3061 0 swss
port 3 n
rlabel metal2 1498 3019 1540 3061 0 b2
port 6 n
rlabel space 1540 3442 1582 3484 0 vctrl
port 7 n
rlabel metal2 2720 -1073 2762 -1031 0 swff
port 1 n
rlabel metal2 1498 -1073 1540 -1031 1 b0
port 4 n
rlabel metal2 1498 973 1540 1015 0 b1
port 5 n
rlabel metal2 2720 973 2762 1015 6 swtt
port 2 n
rlabel metal1 1540 -2564 1582 -2522 4 vctrl
port 8 n
rlabel metal2 2440 -2358 2510 -2288 0 vss
port 9 n
rlabel metal2 1801 -2455 1871 -2385 0 vdd
port 10 n
<< end >>
