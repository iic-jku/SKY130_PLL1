magic
tech sky130A
magscale 1 2
timestamp 1666514521
<< locali >>
rect -81 244 -16 259
rect -81 208 -66 244
rect -30 208 -16 244
rect 274 246 330 261
rect -81 193 -16 208
rect 274 210 284 246
rect 320 210 330 246
rect 1843 256 1909 265
rect 1843 220 1858 256
rect 1894 220 1909 256
rect 1843 211 1909 220
rect 2013 256 2079 265
rect 2013 220 2028 256
rect 2064 220 2079 256
rect 2013 211 2079 220
rect 274 195 330 210
rect 1937 119 1985 125
rect 1937 85 1944 119
rect 1978 85 1985 119
rect 1937 78 1985 85
rect 1380 -129 1446 -114
rect 1380 -165 1395 -129
rect 1431 -165 1446 -129
rect 1421 -180 1446 -165
rect 274 -210 330 -195
rect 274 -246 284 -210
rect 320 -246 330 -210
rect 274 -261 330 -246
rect 274 -842 330 -827
rect 274 -878 284 -842
rect 320 -878 330 -842
rect 274 -893 330 -878
rect 1422 -923 1446 -908
rect 1380 -959 1395 -923
rect 1431 -959 1446 -923
rect 1380 -974 1446 -959
rect 1380 -1217 1446 -1202
rect 1380 -1253 1395 -1217
rect 1431 -1253 1446 -1217
rect 1422 -1268 1446 -1253
rect 16 -1299 82 -1284
rect 16 -1335 31 -1299
rect 67 -1335 82 -1299
rect 16 -1350 82 -1335
rect 274 -1298 330 -1283
rect 274 -1334 284 -1298
rect 320 -1334 330 -1298
rect 274 -1349 330 -1334
rect 1663 -1396 1729 -1387
rect 1663 -1432 1678 -1396
rect 1714 -1432 1729 -1396
rect 1663 -1447 1729 -1432
<< viali >>
rect -66 208 -30 244
rect 29 212 69 252
rect 284 210 320 246
rect 1858 220 1894 256
rect 2028 220 2064 256
rect 1395 129 1431 165
rect 1944 85 1978 119
rect 1395 -165 1431 -129
rect 29 -252 69 -212
rect 284 -246 320 -210
rect 29 -876 69 -836
rect 284 -878 320 -842
rect 1395 -959 1431 -923
rect 1395 -1253 1431 -1217
rect 31 -1335 67 -1299
rect 284 -1334 320 -1298
rect 1678 -1432 1714 -1396
<< metal1 >>
rect 1748 496 1824 592
rect -81 252 -16 259
rect 22 252 78 265
rect 1843 264 1909 271
rect -81 200 -74 252
rect -22 212 29 252
rect 69 212 78 252
rect -22 200 78 212
rect -81 199 78 200
rect 269 254 335 261
rect 269 202 276 254
rect 328 248 335 254
rect 328 208 1528 248
rect 328 202 335 208
rect -81 193 -16 199
rect 269 195 335 202
rect -68 -199 -28 193
rect 1380 173 1446 180
rect 1380 121 1387 173
rect 1439 121 1446 173
rect 1380 114 1446 121
rect 1488 122 1528 208
rect 1843 212 1850 264
rect 1902 212 1909 264
rect 1843 205 1909 212
rect 2013 264 2079 271
rect 2013 212 2020 264
rect 2072 212 2079 264
rect 2013 205 2079 212
rect 1932 122 1990 131
rect 1488 119 1990 122
rect 1488 85 1944 119
rect 1978 85 1990 119
rect 1488 82 1990 85
rect 1932 76 1990 82
rect 1748 -48 1824 48
rect 1380 -121 1446 -114
rect 1380 -173 1387 -121
rect 1439 -127 1446 -121
rect 1844 -127 1850 -121
rect 1439 -167 1850 -127
rect 1439 -173 1446 -167
rect 1844 -173 1850 -167
rect 1902 -173 1908 -121
rect 1380 -180 1446 -173
rect -68 -212 78 -199
rect -68 -252 29 -212
rect 69 -252 78 -212
rect -68 -265 78 -252
rect 269 -202 335 -195
rect 269 -254 276 -202
rect 328 -254 335 -202
rect 269 -261 335 -254
rect -68 -823 -28 -265
rect -68 -836 78 -823
rect -68 -876 29 -836
rect 69 -876 78 -836
rect 22 -889 78 -876
rect 269 -834 335 -827
rect 269 -886 276 -834
rect 328 -886 335 -834
rect 269 -893 335 -886
rect 1380 -915 1446 -908
rect 1380 -967 1387 -915
rect 1439 -921 1446 -915
rect 2013 -921 2019 -915
rect 1439 -961 2019 -921
rect 1439 -967 1446 -961
rect 2013 -967 2019 -961
rect 2071 -967 2077 -915
rect 1380 -974 1446 -967
rect 1380 -1209 1446 -1202
rect 1380 -1261 1387 -1209
rect 1439 -1261 1446 -1209
rect 1380 -1268 1446 -1261
rect 16 -1297 82 -1284
rect 269 -1290 335 -1283
rect 146 -1297 152 -1291
rect 16 -1299 152 -1297
rect 16 -1335 31 -1299
rect 67 -1335 152 -1299
rect 16 -1337 152 -1335
rect 16 -1350 82 -1337
rect 146 -1343 152 -1337
rect 204 -1343 210 -1291
rect 269 -1342 276 -1290
rect 328 -1342 335 -1290
rect 269 -1349 335 -1342
rect 1663 -1388 1729 -1381
rect 1663 -1440 1670 -1388
rect 1722 -1440 1729 -1388
rect 1663 -1447 1729 -1440
<< via1 >>
rect 20 518 72 570
rect -74 244 -22 252
rect -74 208 -66 244
rect -66 208 -30 244
rect -30 208 -22 244
rect -74 200 -22 208
rect 276 246 328 254
rect 276 210 284 246
rect 284 210 320 246
rect 320 210 328 246
rect 276 202 328 210
rect 1387 165 1439 173
rect 1387 129 1395 165
rect 1395 129 1431 165
rect 1431 129 1439 165
rect 1387 121 1439 129
rect 1850 256 1902 264
rect 1850 220 1858 256
rect 1858 220 1894 256
rect 1894 220 1902 256
rect 1850 212 1902 220
rect 2020 256 2072 264
rect 2020 220 2028 256
rect 2028 220 2064 256
rect 2064 220 2072 256
rect 2020 212 2072 220
rect 1676 -26 1728 26
rect 1387 -129 1439 -121
rect 1387 -165 1395 -129
rect 1395 -165 1431 -129
rect 1431 -165 1439 -129
rect 1387 -173 1439 -165
rect 1850 -173 1902 -121
rect 276 -210 328 -202
rect 276 -246 284 -210
rect 284 -246 320 -210
rect 320 -246 328 -210
rect 276 -254 328 -246
rect 20 -570 72 -518
rect 276 -842 328 -834
rect 276 -878 284 -842
rect 284 -878 320 -842
rect 320 -878 328 -842
rect 276 -886 328 -878
rect 1387 -923 1439 -915
rect 1387 -959 1395 -923
rect 1395 -959 1431 -923
rect 1431 -959 1439 -923
rect 1387 -967 1439 -959
rect 2019 -967 2071 -915
rect 1676 -1114 1728 -1062
rect 1387 -1217 1439 -1209
rect 1387 -1253 1395 -1217
rect 1395 -1253 1431 -1217
rect 1431 -1253 1439 -1217
rect 1387 -1261 1439 -1253
rect 152 -1343 204 -1291
rect 276 -1298 328 -1290
rect 276 -1334 284 -1298
rect 284 -1334 320 -1298
rect 320 -1334 328 -1298
rect 276 -1342 328 -1334
rect 1670 -1396 1722 -1388
rect 1670 -1432 1678 -1396
rect 1678 -1432 1714 -1396
rect 1714 -1432 1722 -1396
rect 1670 -1440 1722 -1432
rect 20 -1658 72 -1606
<< metal2 >>
rect 14 570 78 697
rect 14 518 20 570
rect 72 518 78 570
rect -81 252 -16 259
rect -81 200 -74 252
rect -22 200 -16 252
rect -81 193 -16 200
rect 14 -518 78 518
rect 269 254 335 261
rect 269 202 276 254
rect 328 202 335 254
rect 269 195 335 202
rect 1380 173 1446 180
rect 1380 167 1387 173
rect 282 127 1387 167
rect 282 -195 322 127
rect 1380 121 1387 127
rect 1439 121 1446 173
rect 1380 114 1446 121
rect 1670 26 1734 697
rect 1843 264 1909 271
rect 1843 212 1850 264
rect 1902 212 1909 264
rect 1843 205 1909 212
rect 2013 264 2079 271
rect 2013 212 2020 264
rect 2072 212 2079 264
rect 2013 205 2079 212
rect 1670 -26 1676 26
rect 1728 -26 1734 26
rect 1380 -121 1446 -114
rect 1380 -173 1387 -121
rect 1439 -173 1446 -121
rect 1380 -180 1446 -173
rect 269 -202 335 -195
rect 269 -208 276 -202
rect 14 -570 20 -518
rect 72 -570 78 -518
rect 14 -1606 78 -570
rect 158 -248 276 -208
rect 158 -1285 198 -248
rect 269 -254 276 -248
rect 328 -254 335 -202
rect 269 -261 335 -254
rect 269 -834 335 -827
rect 269 -886 276 -834
rect 328 -840 335 -834
rect 1393 -840 1433 -180
rect 328 -880 1433 -840
rect 328 -886 335 -880
rect 269 -893 335 -886
rect 1380 -915 1446 -908
rect 1380 -967 1387 -915
rect 1439 -967 1446 -915
rect 1380 -974 1446 -967
rect 1670 -1062 1734 -26
rect 1856 -115 1896 205
rect 1850 -121 1902 -115
rect 1850 -179 1902 -173
rect 2025 -909 2065 205
rect 2019 -915 2071 -909
rect 2019 -973 2071 -967
rect 1670 -1114 1676 -1062
rect 1728 -1114 1734 -1062
rect 1670 -1121 1734 -1114
rect 1380 -1209 1446 -1202
rect 1380 -1261 1387 -1209
rect 1439 -1215 1446 -1209
rect 1439 -1255 1861 -1215
rect 1439 -1261 1446 -1255
rect 1380 -1268 1446 -1261
rect 152 -1291 204 -1285
rect 152 -1349 204 -1343
rect 269 -1290 335 -1283
rect 269 -1342 276 -1290
rect 328 -1296 335 -1290
rect 328 -1336 1716 -1296
rect 328 -1342 335 -1336
rect 269 -1349 335 -1342
rect 1676 -1381 1716 -1336
rect 1663 -1388 1729 -1381
rect 1663 -1440 1670 -1388
rect 1722 -1440 1729 -1388
rect 1663 -1447 1729 -1440
rect 14 -1658 20 -1606
rect 72 -1658 78 -1606
rect 14 -1665 78 -1658
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 0 0 1 0
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_1
timestamp 1644511149
transform 1 0 0 0 -1 0
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_2
timestamp 1644511149
transform 1 0 0 0 1 -1088
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_3
timestamp 1644511149
transform 1 0 0 0 -1 -1088
box -38 -48 1786 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1824 0 1 0
box -38 -48 314 592
<< labels >>
rlabel metal2 1821 -1255 1861 -1215 0 clk_out
rlabel metal1 -68 -265 -2 -199 0 clk_in
rlabel metal2 14 633 78 697 0 vdd
rlabel metal2 1670 633 1734 697 5 vss
<< end >>
