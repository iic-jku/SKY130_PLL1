magic
tech sky130A
magscale 1 2
timestamp 1668108937
<< metal3 >>
rect -3186 66750 -1463 67041
rect 3185 66750 4908 67041
rect 9556 66750 11279 67041
rect 15927 66750 17650 67041
rect 22298 66750 24021 67041
rect 28669 66750 30392 67041
rect 35040 66750 36763 67041
rect 41411 66750 43134 67041
rect 47782 66750 49505 67041
rect 54153 66750 55876 67041
rect -3186 62393 2894 66750
rect 3185 62393 9265 66750
rect 9556 62393 15636 66750
rect 15927 62393 22007 66750
rect 22298 62393 28378 66750
rect 28669 62393 34749 66750
rect 35040 62393 41120 66750
rect 41411 62393 47491 66750
rect 47782 62393 53862 66750
rect 54153 62393 60233 66750
rect -3186 60670 60524 62393
rect -3186 60379 -1463 60670
rect 3185 60379 4908 60670
rect 9556 60379 11279 60670
rect 15927 60379 17650 60670
rect 22298 60379 24021 60670
rect 28669 60379 30392 60670
rect 35040 60379 36763 60670
rect 41411 60379 43134 60670
rect 47782 60379 49505 60670
rect 54153 60379 55876 60670
rect -3186 56022 2894 60379
rect 3185 56022 9265 60379
rect 9556 56022 15636 60379
rect 15927 56022 22007 60379
rect 22298 56022 28378 60379
rect 28669 56022 34749 60379
rect 35040 56022 41120 60379
rect 41411 56022 47491 60379
rect 47782 56022 53862 60379
rect 54153 56022 60233 60379
rect -3186 54299 60524 56022
rect -3186 54008 -1463 54299
rect 3185 54008 4908 54299
rect 9556 54008 11279 54299
rect 15927 54008 17650 54299
rect 22298 54008 24021 54299
rect 28669 54008 30392 54299
rect 35040 54008 36763 54299
rect 41411 54008 43134 54299
rect 47782 54008 49505 54299
rect 54153 54008 55876 54299
rect -3186 49651 2894 54008
rect 3185 49651 9265 54008
rect 9556 49651 15636 54008
rect 15927 49651 22007 54008
rect 22298 49651 28378 54008
rect 28669 49651 34749 54008
rect 35040 49651 41120 54008
rect 41411 49651 47491 54008
rect 47782 49651 53862 54008
rect 54153 49651 60233 54008
rect -3186 47928 60524 49651
rect -3186 47637 -1463 47928
rect 3185 47637 4908 47928
rect 9556 47637 11279 47928
rect 15927 47637 17650 47928
rect 22298 47637 24021 47928
rect 28669 47637 30392 47928
rect 35040 47637 36763 47928
rect 41411 47637 43134 47928
rect 47782 47637 49505 47928
rect 54153 47637 55876 47928
rect -3186 43280 2894 47637
rect 3185 43280 9265 47637
rect 9556 43280 15636 47637
rect 15927 43280 22007 47637
rect 22298 43280 28378 47637
rect 28669 43280 34749 47637
rect 35040 43280 41120 47637
rect 41411 43280 47491 47637
rect 47782 43280 53862 47637
rect 54153 43280 60233 47637
rect -3186 41557 60524 43280
rect -3186 41266 -1463 41557
rect 3185 41266 4908 41557
rect 9556 41266 11279 41557
rect 15927 41266 17650 41557
rect 22298 41266 24021 41557
rect 28669 41266 30392 41557
rect 35040 41266 36763 41557
rect 41411 41266 43134 41557
rect 47782 41266 49505 41557
rect 54153 41266 55876 41557
rect -3186 36909 2894 41266
rect 3185 36909 9265 41266
rect 9556 36909 15636 41266
rect 15927 36909 22007 41266
rect 22298 36909 28378 41266
rect 28669 36909 34749 41266
rect 35040 36909 41120 41266
rect 41411 36909 47491 41266
rect 47782 36909 53862 41266
rect 54153 36909 60233 41266
rect -3186 35186 60524 36909
rect -3186 34895 -1463 35186
rect 3185 34895 4908 35186
rect 9556 34895 11279 35186
rect 15927 34895 17650 35186
rect 22298 34895 24021 35186
rect 28669 34895 30392 35186
rect 35040 34895 36763 35186
rect 41411 34895 43134 35186
rect 47782 34895 49505 35186
rect 54153 34895 55876 35186
rect -3186 30538 2894 34895
rect 3185 30538 9265 34895
rect 9556 30538 15636 34895
rect 15927 30538 22007 34895
rect 22298 30538 28378 34895
rect 28669 30538 34749 34895
rect 35040 30538 41120 34895
rect 41411 30538 47491 34895
rect 47782 30538 53862 34895
rect 54153 30538 60233 34895
rect -3186 28815 60524 30538
rect -3186 28524 -1463 28815
rect 3185 28524 4908 28815
rect 9556 28524 11279 28815
rect 15927 28524 17650 28815
rect 22298 28524 24021 28815
rect 28669 28524 30392 28815
rect 35040 28524 36763 28815
rect 41411 28524 43134 28815
rect 47782 28524 49505 28815
rect 54153 28524 55876 28815
rect -3186 24167 2894 28524
rect 3185 24167 9265 28524
rect 9556 24167 15636 28524
rect 15927 24167 22007 28524
rect 22298 24167 28378 28524
rect 28669 24167 34749 28524
rect 35040 24167 41120 28524
rect 41411 24167 47491 28524
rect 47782 24167 53862 28524
rect 54153 24167 60233 28524
rect -3186 22444 60524 24167
rect -3186 22153 -1463 22444
rect 3185 22153 4908 22444
rect 9556 22153 11279 22444
rect 15927 22153 17650 22444
rect 22298 22153 24021 22444
rect 28669 22153 30392 22444
rect 35040 22153 36763 22444
rect 41411 22153 43134 22444
rect 47782 22153 49505 22444
rect 54153 22153 55876 22444
rect -3186 17796 2894 22153
rect 3185 17796 9265 22153
rect 9556 17796 15636 22153
rect 15927 17796 22007 22153
rect 22298 17796 28378 22153
rect 28669 17796 34749 22153
rect 35040 17796 41120 22153
rect 41411 17796 47491 22153
rect 47782 17796 53862 22153
rect 54153 17796 60233 22153
rect -3186 16073 60524 17796
rect -3186 15782 -1463 16073
rect 3185 15782 4908 16073
rect 9556 15782 11279 16073
rect 15927 15782 17650 16073
rect 22298 15782 24021 16073
rect 28669 15782 30392 16073
rect 35040 15782 36763 16073
rect 41411 15782 43134 16073
rect 47782 15782 49505 16073
rect 54153 15782 55876 16073
rect -3186 11425 2894 15782
rect 3185 11425 9265 15782
rect 9556 11425 15636 15782
rect 15927 11425 22007 15782
rect 22298 11425 28378 15782
rect 28669 11425 34749 15782
rect 35040 11425 41120 15782
rect 41411 11425 47491 15782
rect 47782 11425 53862 15782
rect 54153 11425 60233 15782
rect -3186 9702 60524 11425
rect -3186 9411 -1463 9702
rect 3185 9411 4908 9702
rect 9556 9411 11279 9702
rect 15927 9411 17650 9702
rect 22298 9411 24021 9702
rect 28669 9411 30392 9702
rect 35040 9411 36763 9702
rect 41411 9411 43134 9702
rect 47782 9411 49505 9702
rect 54153 9411 55876 9702
rect -3186 5054 2894 9411
rect 3185 5054 9265 9411
rect 9556 5054 15636 9411
rect 15927 5054 22007 9411
rect 22298 5054 28378 9411
rect 28669 5054 34749 9411
rect 35040 5054 41120 9411
rect 41411 5054 47491 9411
rect 47782 5054 53862 9411
rect 54153 5054 60233 9411
rect -3186 3331 60524 5054
rect -3186 3040 -1463 3331
rect 3185 3040 4908 3331
rect 9556 3040 11279 3331
rect 15927 3040 17650 3331
rect 22298 3040 24021 3331
rect 28669 3040 30392 3331
rect 35040 3040 36763 3331
rect 41411 3040 43134 3331
rect 47782 3040 49505 3331
rect 54153 3040 55876 3331
rect -3186 -1317 2894 3040
rect 3185 -1317 9265 3040
rect 9556 -1317 15636 3040
rect 15927 -1317 22007 3040
rect 22298 -1317 28378 3040
rect 28669 -1317 34749 3040
rect 35040 -1317 41120 3040
rect 41411 -1317 47491 3040
rect 47782 -1317 53862 3040
rect 54153 -1317 60233 3040
rect -3186 -3040 60524 -1317
<< mimcap >>
rect -3146 66670 2854 66710
rect -3146 60750 -3106 66670
rect 2814 60750 2854 66670
rect -3146 60710 2854 60750
rect 3225 66670 9225 66710
rect 3225 60750 3265 66670
rect 9185 60750 9225 66670
rect 3225 60710 9225 60750
rect 9596 66670 15596 66710
rect 9596 60750 9636 66670
rect 15556 60750 15596 66670
rect 9596 60710 15596 60750
rect 15967 66670 21967 66710
rect 15967 60750 16007 66670
rect 21927 60750 21967 66670
rect 15967 60710 21967 60750
rect 22338 66670 28338 66710
rect 22338 60750 22378 66670
rect 28298 60750 28338 66670
rect 22338 60710 28338 60750
rect 28709 66670 34709 66710
rect 28709 60750 28749 66670
rect 34669 60750 34709 66670
rect 28709 60710 34709 60750
rect 35080 66670 41080 66710
rect 35080 60750 35120 66670
rect 41040 60750 41080 66670
rect 35080 60710 41080 60750
rect 41451 66670 47451 66710
rect 41451 60750 41491 66670
rect 47411 60750 47451 66670
rect 41451 60710 47451 60750
rect 47822 66670 53822 66710
rect 47822 60750 47862 66670
rect 53782 60750 53822 66670
rect 47822 60710 53822 60750
rect 54193 66670 60193 66710
rect 54193 60750 54233 66670
rect 60153 60750 60193 66670
rect 54193 60710 60193 60750
rect -3146 60299 2854 60339
rect -3146 54379 -3106 60299
rect 2814 54379 2854 60299
rect -3146 54339 2854 54379
rect 3225 60299 9225 60339
rect 3225 54379 3265 60299
rect 9185 54379 9225 60299
rect 3225 54339 9225 54379
rect 9596 60299 15596 60339
rect 9596 54379 9636 60299
rect 15556 54379 15596 60299
rect 9596 54339 15596 54379
rect 15967 60299 21967 60339
rect 15967 54379 16007 60299
rect 21927 54379 21967 60299
rect 15967 54339 21967 54379
rect 22338 60299 28338 60339
rect 22338 54379 22378 60299
rect 28298 54379 28338 60299
rect 22338 54339 28338 54379
rect 28709 60299 34709 60339
rect 28709 54379 28749 60299
rect 34669 54379 34709 60299
rect 28709 54339 34709 54379
rect 35080 60299 41080 60339
rect 35080 54379 35120 60299
rect 41040 54379 41080 60299
rect 35080 54339 41080 54379
rect 41451 60299 47451 60339
rect 41451 54379 41491 60299
rect 47411 54379 47451 60299
rect 41451 54339 47451 54379
rect 47822 60299 53822 60339
rect 47822 54379 47862 60299
rect 53782 54379 53822 60299
rect 47822 54339 53822 54379
rect 54193 60299 60193 60339
rect 54193 54379 54233 60299
rect 60153 54379 60193 60299
rect 54193 54339 60193 54379
rect -3146 53928 2854 53968
rect -3146 48008 -3106 53928
rect 2814 48008 2854 53928
rect -3146 47968 2854 48008
rect 3225 53928 9225 53968
rect 3225 48008 3265 53928
rect 9185 48008 9225 53928
rect 3225 47968 9225 48008
rect 9596 53928 15596 53968
rect 9596 48008 9636 53928
rect 15556 48008 15596 53928
rect 9596 47968 15596 48008
rect 15967 53928 21967 53968
rect 15967 48008 16007 53928
rect 21927 48008 21967 53928
rect 15967 47968 21967 48008
rect 22338 53928 28338 53968
rect 22338 48008 22378 53928
rect 28298 48008 28338 53928
rect 22338 47968 28338 48008
rect 28709 53928 34709 53968
rect 28709 48008 28749 53928
rect 34669 48008 34709 53928
rect 28709 47968 34709 48008
rect 35080 53928 41080 53968
rect 35080 48008 35120 53928
rect 41040 48008 41080 53928
rect 35080 47968 41080 48008
rect 41451 53928 47451 53968
rect 41451 48008 41491 53928
rect 47411 48008 47451 53928
rect 41451 47968 47451 48008
rect 47822 53928 53822 53968
rect 47822 48008 47862 53928
rect 53782 48008 53822 53928
rect 47822 47968 53822 48008
rect 54193 53928 60193 53968
rect 54193 48008 54233 53928
rect 60153 48008 60193 53928
rect 54193 47968 60193 48008
rect -3146 47557 2854 47597
rect -3146 41637 -3106 47557
rect 2814 41637 2854 47557
rect -3146 41597 2854 41637
rect 3225 47557 9225 47597
rect 3225 41637 3265 47557
rect 9185 41637 9225 47557
rect 3225 41597 9225 41637
rect 9596 47557 15596 47597
rect 9596 41637 9636 47557
rect 15556 41637 15596 47557
rect 9596 41597 15596 41637
rect 15967 47557 21967 47597
rect 15967 41637 16007 47557
rect 21927 41637 21967 47557
rect 15967 41597 21967 41637
rect 22338 47557 28338 47597
rect 22338 41637 22378 47557
rect 28298 41637 28338 47557
rect 22338 41597 28338 41637
rect 28709 47557 34709 47597
rect 28709 41637 28749 47557
rect 34669 41637 34709 47557
rect 28709 41597 34709 41637
rect 35080 47557 41080 47597
rect 35080 41637 35120 47557
rect 41040 41637 41080 47557
rect 35080 41597 41080 41637
rect 41451 47557 47451 47597
rect 41451 41637 41491 47557
rect 47411 41637 47451 47557
rect 41451 41597 47451 41637
rect 47822 47557 53822 47597
rect 47822 41637 47862 47557
rect 53782 41637 53822 47557
rect 47822 41597 53822 41637
rect 54193 47557 60193 47597
rect 54193 41637 54233 47557
rect 60153 41637 60193 47557
rect 54193 41597 60193 41637
rect -3146 41186 2854 41226
rect -3146 35266 -3106 41186
rect 2814 35266 2854 41186
rect -3146 35226 2854 35266
rect 3225 41186 9225 41226
rect 3225 35266 3265 41186
rect 9185 35266 9225 41186
rect 3225 35226 9225 35266
rect 9596 41186 15596 41226
rect 9596 35266 9636 41186
rect 15556 35266 15596 41186
rect 9596 35226 15596 35266
rect 15967 41186 21967 41226
rect 15967 35266 16007 41186
rect 21927 35266 21967 41186
rect 15967 35226 21967 35266
rect 22338 41186 28338 41226
rect 22338 35266 22378 41186
rect 28298 35266 28338 41186
rect 22338 35226 28338 35266
rect 28709 41186 34709 41226
rect 28709 35266 28749 41186
rect 34669 35266 34709 41186
rect 28709 35226 34709 35266
rect 35080 41186 41080 41226
rect 35080 35266 35120 41186
rect 41040 35266 41080 41186
rect 35080 35226 41080 35266
rect 41451 41186 47451 41226
rect 41451 35266 41491 41186
rect 47411 35266 47451 41186
rect 41451 35226 47451 35266
rect 47822 41186 53822 41226
rect 47822 35266 47862 41186
rect 53782 35266 53822 41186
rect 47822 35226 53822 35266
rect 54193 41186 60193 41226
rect 54193 35266 54233 41186
rect 60153 35266 60193 41186
rect 54193 35226 60193 35266
rect -3146 34815 2854 34855
rect -3146 28895 -3106 34815
rect 2814 28895 2854 34815
rect -3146 28855 2854 28895
rect 3225 34815 9225 34855
rect 3225 28895 3265 34815
rect 9185 28895 9225 34815
rect 3225 28855 9225 28895
rect 9596 34815 15596 34855
rect 9596 28895 9636 34815
rect 15556 28895 15596 34815
rect 9596 28855 15596 28895
rect 15967 34815 21967 34855
rect 15967 28895 16007 34815
rect 21927 28895 21967 34815
rect 15967 28855 21967 28895
rect 22338 34815 28338 34855
rect 22338 28895 22378 34815
rect 28298 28895 28338 34815
rect 22338 28855 28338 28895
rect 28709 34815 34709 34855
rect 28709 28895 28749 34815
rect 34669 28895 34709 34815
rect 28709 28855 34709 28895
rect 35080 34815 41080 34855
rect 35080 28895 35120 34815
rect 41040 28895 41080 34815
rect 35080 28855 41080 28895
rect 41451 34815 47451 34855
rect 41451 28895 41491 34815
rect 47411 28895 47451 34815
rect 41451 28855 47451 28895
rect 47822 34815 53822 34855
rect 47822 28895 47862 34815
rect 53782 28895 53822 34815
rect 47822 28855 53822 28895
rect 54193 34815 60193 34855
rect 54193 28895 54233 34815
rect 60153 28895 60193 34815
rect 54193 28855 60193 28895
rect -3146 28444 2854 28484
rect -3146 22524 -3106 28444
rect 2814 22524 2854 28444
rect -3146 22484 2854 22524
rect 3225 28444 9225 28484
rect 3225 22524 3265 28444
rect 9185 22524 9225 28444
rect 3225 22484 9225 22524
rect 9596 28444 15596 28484
rect 9596 22524 9636 28444
rect 15556 22524 15596 28444
rect 9596 22484 15596 22524
rect 15967 28444 21967 28484
rect 15967 22524 16007 28444
rect 21927 22524 21967 28444
rect 15967 22484 21967 22524
rect 22338 28444 28338 28484
rect 22338 22524 22378 28444
rect 28298 22524 28338 28444
rect 22338 22484 28338 22524
rect 28709 28444 34709 28484
rect 28709 22524 28749 28444
rect 34669 22524 34709 28444
rect 28709 22484 34709 22524
rect 35080 28444 41080 28484
rect 35080 22524 35120 28444
rect 41040 22524 41080 28444
rect 35080 22484 41080 22524
rect 41451 28444 47451 28484
rect 41451 22524 41491 28444
rect 47411 22524 47451 28444
rect 41451 22484 47451 22524
rect 47822 28444 53822 28484
rect 47822 22524 47862 28444
rect 53782 22524 53822 28444
rect 47822 22484 53822 22524
rect 54193 28444 60193 28484
rect 54193 22524 54233 28444
rect 60153 22524 60193 28444
rect 54193 22484 60193 22524
rect -3146 22073 2854 22113
rect -3146 16153 -3106 22073
rect 2814 16153 2854 22073
rect -3146 16113 2854 16153
rect 3225 22073 9225 22113
rect 3225 16153 3265 22073
rect 9185 16153 9225 22073
rect 3225 16113 9225 16153
rect 9596 22073 15596 22113
rect 9596 16153 9636 22073
rect 15556 16153 15596 22073
rect 9596 16113 15596 16153
rect 15967 22073 21967 22113
rect 15967 16153 16007 22073
rect 21927 16153 21967 22073
rect 15967 16113 21967 16153
rect 22338 22073 28338 22113
rect 22338 16153 22378 22073
rect 28298 16153 28338 22073
rect 22338 16113 28338 16153
rect 28709 22073 34709 22113
rect 28709 16153 28749 22073
rect 34669 16153 34709 22073
rect 28709 16113 34709 16153
rect 35080 22073 41080 22113
rect 35080 16153 35120 22073
rect 41040 16153 41080 22073
rect 35080 16113 41080 16153
rect 41451 22073 47451 22113
rect 41451 16153 41491 22073
rect 47411 16153 47451 22073
rect 41451 16113 47451 16153
rect 47822 22073 53822 22113
rect 47822 16153 47862 22073
rect 53782 16153 53822 22073
rect 47822 16113 53822 16153
rect 54193 22073 60193 22113
rect 54193 16153 54233 22073
rect 60153 16153 60193 22073
rect 54193 16113 60193 16153
rect -3146 15702 2854 15742
rect -3146 9782 -3106 15702
rect 2814 9782 2854 15702
rect -3146 9742 2854 9782
rect 3225 15702 9225 15742
rect 3225 9782 3265 15702
rect 9185 9782 9225 15702
rect 3225 9742 9225 9782
rect 9596 15702 15596 15742
rect 9596 9782 9636 15702
rect 15556 9782 15596 15702
rect 9596 9742 15596 9782
rect 15967 15702 21967 15742
rect 15967 9782 16007 15702
rect 21927 9782 21967 15702
rect 15967 9742 21967 9782
rect 22338 15702 28338 15742
rect 22338 9782 22378 15702
rect 28298 9782 28338 15702
rect 22338 9742 28338 9782
rect 28709 15702 34709 15742
rect 28709 9782 28749 15702
rect 34669 9782 34709 15702
rect 28709 9742 34709 9782
rect 35080 15702 41080 15742
rect 35080 9782 35120 15702
rect 41040 9782 41080 15702
rect 35080 9742 41080 9782
rect 41451 15702 47451 15742
rect 41451 9782 41491 15702
rect 47411 9782 47451 15702
rect 41451 9742 47451 9782
rect 47822 15702 53822 15742
rect 47822 9782 47862 15702
rect 53782 9782 53822 15702
rect 47822 9742 53822 9782
rect 54193 15702 60193 15742
rect 54193 9782 54233 15702
rect 60153 9782 60193 15702
rect 54193 9742 60193 9782
rect -3146 9331 2854 9371
rect -3146 3411 -3106 9331
rect 2814 3411 2854 9331
rect -3146 3371 2854 3411
rect 3225 9331 9225 9371
rect 3225 3411 3265 9331
rect 9185 3411 9225 9331
rect 3225 3371 9225 3411
rect 9596 9331 15596 9371
rect 9596 3411 9636 9331
rect 15556 3411 15596 9331
rect 9596 3371 15596 3411
rect 15967 9331 21967 9371
rect 15967 3411 16007 9331
rect 21927 3411 21967 9331
rect 15967 3371 21967 3411
rect 22338 9331 28338 9371
rect 22338 3411 22378 9331
rect 28298 3411 28338 9331
rect 22338 3371 28338 3411
rect 28709 9331 34709 9371
rect 28709 3411 28749 9331
rect 34669 3411 34709 9331
rect 28709 3371 34709 3411
rect 35080 9331 41080 9371
rect 35080 3411 35120 9331
rect 41040 3411 41080 9331
rect 35080 3371 41080 3411
rect 41451 9331 47451 9371
rect 41451 3411 41491 9331
rect 47411 3411 47451 9331
rect 41451 3371 47451 3411
rect 47822 9331 53822 9371
rect 47822 3411 47862 9331
rect 53782 3411 53822 9331
rect 47822 3371 53822 3411
rect 54193 9331 60193 9371
rect 54193 3411 54233 9331
rect 60153 3411 60193 9331
rect 54193 3371 60193 3411
rect -3146 2960 2854 3000
rect -3146 -2960 -3106 2960
rect 2814 -2960 2854 2960
rect -3146 -3000 2854 -2960
rect 3225 2960 9225 3000
rect 3225 -2960 3265 2960
rect 9185 -2960 9225 2960
rect 3225 -3000 9225 -2960
rect 9596 2960 15596 3000
rect 9596 -2960 9636 2960
rect 15556 -2960 15596 2960
rect 9596 -3000 15596 -2960
rect 15967 2960 21967 3000
rect 15967 -2960 16007 2960
rect 21927 -2960 21967 2960
rect 15967 -3000 21967 -2960
rect 22338 2960 28338 3000
rect 22338 -2960 22378 2960
rect 28298 -2960 28338 2960
rect 22338 -3000 28338 -2960
rect 28709 2960 34709 3000
rect 28709 -2960 28749 2960
rect 34669 -2960 34709 2960
rect 28709 -3000 34709 -2960
rect 35080 2960 41080 3000
rect 35080 -2960 35120 2960
rect 41040 -2960 41080 2960
rect 35080 -3000 41080 -2960
rect 41451 2960 47451 3000
rect 41451 -2960 41491 2960
rect 47411 -2960 47451 2960
rect 41451 -3000 47451 -2960
rect 47822 2960 53822 3000
rect 47822 -2960 47862 2960
rect 53782 -2960 53822 2960
rect 47822 -3000 53822 -2960
rect 54193 2960 60193 3000
rect 54193 -2960 54233 2960
rect 60153 -2960 60193 2960
rect 54193 -3000 60193 -2960
<< mimcapcontact >>
rect -3106 60750 2814 66670
rect 3265 60750 9185 66670
rect 9636 60750 15556 66670
rect 16007 60750 21927 66670
rect 22378 60750 28298 66670
rect 28749 60750 34669 66670
rect 35120 60750 41040 66670
rect 41491 60750 47411 66670
rect 47862 60750 53782 66670
rect 54233 60750 60153 66670
rect -3106 54379 2814 60299
rect 3265 54379 9185 60299
rect 9636 54379 15556 60299
rect 16007 54379 21927 60299
rect 22378 54379 28298 60299
rect 28749 54379 34669 60299
rect 35120 54379 41040 60299
rect 41491 54379 47411 60299
rect 47862 54379 53782 60299
rect 54233 54379 60153 60299
rect -3106 48008 2814 53928
rect 3265 48008 9185 53928
rect 9636 48008 15556 53928
rect 16007 48008 21927 53928
rect 22378 48008 28298 53928
rect 28749 48008 34669 53928
rect 35120 48008 41040 53928
rect 41491 48008 47411 53928
rect 47862 48008 53782 53928
rect 54233 48008 60153 53928
rect -3106 41637 2814 47557
rect 3265 41637 9185 47557
rect 9636 41637 15556 47557
rect 16007 41637 21927 47557
rect 22378 41637 28298 47557
rect 28749 41637 34669 47557
rect 35120 41637 41040 47557
rect 41491 41637 47411 47557
rect 47862 41637 53782 47557
rect 54233 41637 60153 47557
rect -3106 35266 2814 41186
rect 3265 35266 9185 41186
rect 9636 35266 15556 41186
rect 16007 35266 21927 41186
rect 22378 35266 28298 41186
rect 28749 35266 34669 41186
rect 35120 35266 41040 41186
rect 41491 35266 47411 41186
rect 47862 35266 53782 41186
rect 54233 35266 60153 41186
rect -3106 28895 2814 34815
rect 3265 28895 9185 34815
rect 9636 28895 15556 34815
rect 16007 28895 21927 34815
rect 22378 28895 28298 34815
rect 28749 28895 34669 34815
rect 35120 28895 41040 34815
rect 41491 28895 47411 34815
rect 47862 28895 53782 34815
rect 54233 28895 60153 34815
rect -3106 22524 2814 28444
rect 3265 22524 9185 28444
rect 9636 22524 15556 28444
rect 16007 22524 21927 28444
rect 22378 22524 28298 28444
rect 28749 22524 34669 28444
rect 35120 22524 41040 28444
rect 41491 22524 47411 28444
rect 47862 22524 53782 28444
rect 54233 22524 60153 28444
rect -3106 16153 2814 22073
rect 3265 16153 9185 22073
rect 9636 16153 15556 22073
rect 16007 16153 21927 22073
rect 22378 16153 28298 22073
rect 28749 16153 34669 22073
rect 35120 16153 41040 22073
rect 41491 16153 47411 22073
rect 47862 16153 53782 22073
rect 54233 16153 60153 22073
rect -3106 9782 2814 15702
rect 3265 9782 9185 15702
rect 9636 9782 15556 15702
rect 16007 9782 21927 15702
rect 22378 9782 28298 15702
rect 28749 9782 34669 15702
rect 35120 9782 41040 15702
rect 41491 9782 47411 15702
rect 47862 9782 53782 15702
rect 54233 9782 60153 15702
rect -3106 3411 2814 9331
rect 3265 3411 9185 9331
rect 9636 3411 15556 9331
rect 16007 3411 21927 9331
rect 22378 3411 28298 9331
rect 28749 3411 34669 9331
rect 35120 3411 41040 9331
rect 41491 3411 47411 9331
rect 47862 3411 53782 9331
rect 54233 3411 60153 9331
rect -3106 -2960 2814 2960
rect 3265 -2960 9185 2960
rect 9636 -2960 15556 2960
rect 16007 -2960 21927 2960
rect 22378 -2960 28298 2960
rect 28749 -2960 34669 2960
rect 35120 -2960 41040 2960
rect 41491 -2960 47411 2960
rect 47862 -2960 53782 2960
rect 54233 -2960 60153 2960
<< metal4 >>
rect -3146 66710 -1463 67041
rect 3225 66710 4908 67041
rect 9596 66710 11279 67041
rect 15967 66710 17650 67041
rect 22338 66710 24021 67041
rect 28709 66710 30392 67041
rect 35080 66710 36763 67041
rect 41451 66710 43134 67041
rect 47822 66710 49505 67041
rect 54193 66710 55876 67041
rect -3146 66670 2854 66710
rect -3146 62393 -3106 66670
rect -3186 60750 -3106 62393
rect 2814 62393 2854 66670
rect 3225 66670 9225 66710
rect 3225 62393 3265 66670
rect 2814 60750 3265 62393
rect 9185 62393 9225 66670
rect 9596 66670 15596 66710
rect 9596 62393 9636 66670
rect 9185 60750 9636 62393
rect 15556 62393 15596 66670
rect 15967 66670 21967 66710
rect 15967 62393 16007 66670
rect 15556 60750 16007 62393
rect 21927 62393 21967 66670
rect 22338 66670 28338 66710
rect 22338 62393 22378 66670
rect 21927 60750 22378 62393
rect 28298 62393 28338 66670
rect 28709 66670 34709 66710
rect 28709 62393 28749 66670
rect 28298 60750 28749 62393
rect 34669 62393 34709 66670
rect 35080 66670 41080 66710
rect 35080 62393 35120 66670
rect 34669 60750 35120 62393
rect 41040 62393 41080 66670
rect 41451 66670 47451 66710
rect 41451 62393 41491 66670
rect 41040 60750 41491 62393
rect 47411 62393 47451 66670
rect 47822 66670 53822 66710
rect 47822 62393 47862 66670
rect 47411 60750 47862 62393
rect 53782 62393 53822 66670
rect 54193 66670 60193 66710
rect 54193 62393 54233 66670
rect 53782 60750 54233 62393
rect 60153 62393 60193 66670
rect 60153 60750 60524 62393
rect -3186 60710 60524 60750
rect -3146 60339 -1463 60710
rect 3225 60339 4908 60710
rect 9596 60339 11279 60710
rect 15967 60339 17650 60710
rect 22338 60339 24021 60710
rect 28709 60339 30392 60710
rect 35080 60339 36763 60710
rect 41451 60339 43134 60710
rect 47822 60339 49505 60710
rect 54193 60339 55876 60710
rect -3146 60299 2854 60339
rect -3146 56022 -3106 60299
rect -3186 54379 -3106 56022
rect 2814 56022 2854 60299
rect 3225 60299 9225 60339
rect 3225 56022 3265 60299
rect 2814 54379 3265 56022
rect 9185 56022 9225 60299
rect 9596 60299 15596 60339
rect 9596 56022 9636 60299
rect 9185 54379 9636 56022
rect 15556 56022 15596 60299
rect 15967 60299 21967 60339
rect 15967 56022 16007 60299
rect 15556 54379 16007 56022
rect 21927 56022 21967 60299
rect 22338 60299 28338 60339
rect 22338 56022 22378 60299
rect 21927 54379 22378 56022
rect 28298 56022 28338 60299
rect 28709 60299 34709 60339
rect 28709 56022 28749 60299
rect 28298 54379 28749 56022
rect 34669 56022 34709 60299
rect 35080 60299 41080 60339
rect 35080 56022 35120 60299
rect 34669 54379 35120 56022
rect 41040 56022 41080 60299
rect 41451 60299 47451 60339
rect 41451 56022 41491 60299
rect 41040 54379 41491 56022
rect 47411 56022 47451 60299
rect 47822 60299 53822 60339
rect 47822 56022 47862 60299
rect 47411 54379 47862 56022
rect 53782 56022 53822 60299
rect 54193 60299 60193 60339
rect 54193 56022 54233 60299
rect 53782 54379 54233 56022
rect 60153 56022 60193 60299
rect 60153 54379 60524 56022
rect -3186 54339 60524 54379
rect -3146 53968 -1463 54339
rect 3225 53968 4908 54339
rect 9596 53968 11279 54339
rect 15967 53968 17650 54339
rect 22338 53968 24021 54339
rect 28709 53968 30392 54339
rect 35080 53968 36763 54339
rect 41451 53968 43134 54339
rect 47822 53968 49505 54339
rect 54193 53968 55876 54339
rect -3146 53928 2854 53968
rect -3146 49651 -3106 53928
rect -3186 48008 -3106 49651
rect 2814 49651 2854 53928
rect 3225 53928 9225 53968
rect 3225 49651 3265 53928
rect 2814 48008 3265 49651
rect 9185 49651 9225 53928
rect 9596 53928 15596 53968
rect 9596 49651 9636 53928
rect 9185 48008 9636 49651
rect 15556 49651 15596 53928
rect 15967 53928 21967 53968
rect 15967 49651 16007 53928
rect 15556 48008 16007 49651
rect 21927 49651 21967 53928
rect 22338 53928 28338 53968
rect 22338 49651 22378 53928
rect 21927 48008 22378 49651
rect 28298 49651 28338 53928
rect 28709 53928 34709 53968
rect 28709 49651 28749 53928
rect 28298 48008 28749 49651
rect 34669 49651 34709 53928
rect 35080 53928 41080 53968
rect 35080 49651 35120 53928
rect 34669 48008 35120 49651
rect 41040 49651 41080 53928
rect 41451 53928 47451 53968
rect 41451 49651 41491 53928
rect 41040 48008 41491 49651
rect 47411 49651 47451 53928
rect 47822 53928 53822 53968
rect 47822 49651 47862 53928
rect 47411 48008 47862 49651
rect 53782 49651 53822 53928
rect 54193 53928 60193 53968
rect 54193 49651 54233 53928
rect 53782 48008 54233 49651
rect 60153 49651 60193 53928
rect 60153 48008 60524 49651
rect -3186 47968 60524 48008
rect -3146 47597 -1463 47968
rect 3225 47597 4908 47968
rect 9596 47597 11279 47968
rect 15967 47597 17650 47968
rect 22338 47597 24021 47968
rect 28709 47597 30392 47968
rect 35080 47597 36763 47968
rect 41451 47597 43134 47968
rect 47822 47597 49505 47968
rect 54193 47597 55876 47968
rect -3146 47557 2854 47597
rect -3146 43280 -3106 47557
rect -3186 41637 -3106 43280
rect 2814 43280 2854 47557
rect 3225 47557 9225 47597
rect 3225 43280 3265 47557
rect 2814 41637 3265 43280
rect 9185 43280 9225 47557
rect 9596 47557 15596 47597
rect 9596 43280 9636 47557
rect 9185 41637 9636 43280
rect 15556 43280 15596 47557
rect 15967 47557 21967 47597
rect 15967 43280 16007 47557
rect 15556 41637 16007 43280
rect 21927 43280 21967 47557
rect 22338 47557 28338 47597
rect 22338 43280 22378 47557
rect 21927 41637 22378 43280
rect 28298 43280 28338 47557
rect 28709 47557 34709 47597
rect 28709 43280 28749 47557
rect 28298 41637 28749 43280
rect 34669 43280 34709 47557
rect 35080 47557 41080 47597
rect 35080 43280 35120 47557
rect 34669 41637 35120 43280
rect 41040 43280 41080 47557
rect 41451 47557 47451 47597
rect 41451 43280 41491 47557
rect 41040 41637 41491 43280
rect 47411 43280 47451 47557
rect 47822 47557 53822 47597
rect 47822 43280 47862 47557
rect 47411 41637 47862 43280
rect 53782 43280 53822 47557
rect 54193 47557 60193 47597
rect 54193 43280 54233 47557
rect 53782 41637 54233 43280
rect 60153 43280 60193 47557
rect 60153 41637 60524 43280
rect -3186 41597 60524 41637
rect -3146 41226 -1463 41597
rect 3225 41226 4908 41597
rect 9596 41226 11279 41597
rect 15967 41226 17650 41597
rect 22338 41226 24021 41597
rect 28709 41226 30392 41597
rect 35080 41226 36763 41597
rect 41451 41226 43134 41597
rect 47822 41226 49505 41597
rect 54193 41226 55876 41597
rect -3146 41186 2854 41226
rect -3146 36909 -3106 41186
rect -3186 35266 -3106 36909
rect 2814 36909 2854 41186
rect 3225 41186 9225 41226
rect 3225 36909 3265 41186
rect 2814 35266 3265 36909
rect 9185 36909 9225 41186
rect 9596 41186 15596 41226
rect 9596 36909 9636 41186
rect 9185 35266 9636 36909
rect 15556 36909 15596 41186
rect 15967 41186 21967 41226
rect 15967 36909 16007 41186
rect 15556 35266 16007 36909
rect 21927 36909 21967 41186
rect 22338 41186 28338 41226
rect 22338 36909 22378 41186
rect 21927 35266 22378 36909
rect 28298 36909 28338 41186
rect 28709 41186 34709 41226
rect 28709 36909 28749 41186
rect 28298 35266 28749 36909
rect 34669 36909 34709 41186
rect 35080 41186 41080 41226
rect 35080 36909 35120 41186
rect 34669 35266 35120 36909
rect 41040 36909 41080 41186
rect 41451 41186 47451 41226
rect 41451 36909 41491 41186
rect 41040 35266 41491 36909
rect 47411 36909 47451 41186
rect 47822 41186 53822 41226
rect 47822 36909 47862 41186
rect 47411 35266 47862 36909
rect 53782 36909 53822 41186
rect 54193 41186 60193 41226
rect 54193 36909 54233 41186
rect 53782 35266 54233 36909
rect 60153 36909 60193 41186
rect 60153 35266 60524 36909
rect -3186 35226 60524 35266
rect -3146 34855 -1463 35226
rect 3225 34855 4908 35226
rect 9596 34855 11279 35226
rect 15967 34855 17650 35226
rect 22338 34855 24021 35226
rect 28709 34855 30392 35226
rect 35080 34855 36763 35226
rect 41451 34855 43134 35226
rect 47822 34855 49505 35226
rect 54193 34855 55876 35226
rect -3146 34815 2854 34855
rect -3146 30538 -3106 34815
rect -3186 28895 -3106 30538
rect 2814 30538 2854 34815
rect 3225 34815 9225 34855
rect 3225 30538 3265 34815
rect 2814 28895 3265 30538
rect 9185 30538 9225 34815
rect 9596 34815 15596 34855
rect 9596 30538 9636 34815
rect 9185 28895 9636 30538
rect 15556 30538 15596 34815
rect 15967 34815 21967 34855
rect 15967 30538 16007 34815
rect 15556 28895 16007 30538
rect 21927 30538 21967 34815
rect 22338 34815 28338 34855
rect 22338 30538 22378 34815
rect 21927 28895 22378 30538
rect 28298 30538 28338 34815
rect 28709 34815 34709 34855
rect 28709 30538 28749 34815
rect 28298 28895 28749 30538
rect 34669 30538 34709 34815
rect 35080 34815 41080 34855
rect 35080 30538 35120 34815
rect 34669 28895 35120 30538
rect 41040 30538 41080 34815
rect 41451 34815 47451 34855
rect 41451 30538 41491 34815
rect 41040 28895 41491 30538
rect 47411 30538 47451 34815
rect 47822 34815 53822 34855
rect 47822 30538 47862 34815
rect 47411 28895 47862 30538
rect 53782 30538 53822 34815
rect 54193 34815 60193 34855
rect 54193 30538 54233 34815
rect 53782 28895 54233 30538
rect 60153 30538 60193 34815
rect 60153 28895 60524 30538
rect -3186 28855 60524 28895
rect -3146 28484 -1463 28855
rect 3225 28484 4908 28855
rect 9596 28484 11279 28855
rect 15967 28484 17650 28855
rect 22338 28484 24021 28855
rect 28709 28484 30392 28855
rect 35080 28484 36763 28855
rect 41451 28484 43134 28855
rect 47822 28484 49505 28855
rect 54193 28484 55876 28855
rect -3146 28444 2854 28484
rect -3146 24167 -3106 28444
rect -3186 22524 -3106 24167
rect 2814 24167 2854 28444
rect 3225 28444 9225 28484
rect 3225 24167 3265 28444
rect 2814 22524 3265 24167
rect 9185 24167 9225 28444
rect 9596 28444 15596 28484
rect 9596 24167 9636 28444
rect 9185 22524 9636 24167
rect 15556 24167 15596 28444
rect 15967 28444 21967 28484
rect 15967 24167 16007 28444
rect 15556 22524 16007 24167
rect 21927 24167 21967 28444
rect 22338 28444 28338 28484
rect 22338 24167 22378 28444
rect 21927 22524 22378 24167
rect 28298 24167 28338 28444
rect 28709 28444 34709 28484
rect 28709 24167 28749 28444
rect 28298 22524 28749 24167
rect 34669 24167 34709 28444
rect 35080 28444 41080 28484
rect 35080 24167 35120 28444
rect 34669 22524 35120 24167
rect 41040 24167 41080 28444
rect 41451 28444 47451 28484
rect 41451 24167 41491 28444
rect 41040 22524 41491 24167
rect 47411 24167 47451 28444
rect 47822 28444 53822 28484
rect 47822 24167 47862 28444
rect 47411 22524 47862 24167
rect 53782 24167 53822 28444
rect 54193 28444 60193 28484
rect 54193 24167 54233 28444
rect 53782 22524 54233 24167
rect 60153 24167 60193 28444
rect 60153 22524 60524 24167
rect -3186 22484 60524 22524
rect -3146 22113 -1463 22484
rect 3225 22113 4908 22484
rect 9596 22113 11279 22484
rect 15967 22113 17650 22484
rect 22338 22113 24021 22484
rect 28709 22113 30392 22484
rect 35080 22113 36763 22484
rect 41451 22113 43134 22484
rect 47822 22113 49505 22484
rect 54193 22113 55876 22484
rect -3146 22073 2854 22113
rect -3146 17796 -3106 22073
rect -3186 16153 -3106 17796
rect 2814 17796 2854 22073
rect 3225 22073 9225 22113
rect 3225 17796 3265 22073
rect 2814 16153 3265 17796
rect 9185 17796 9225 22073
rect 9596 22073 15596 22113
rect 9596 17796 9636 22073
rect 9185 16153 9636 17796
rect 15556 17796 15596 22073
rect 15967 22073 21967 22113
rect 15967 17796 16007 22073
rect 15556 16153 16007 17796
rect 21927 17796 21967 22073
rect 22338 22073 28338 22113
rect 22338 17796 22378 22073
rect 21927 16153 22378 17796
rect 28298 17796 28338 22073
rect 28709 22073 34709 22113
rect 28709 17796 28749 22073
rect 28298 16153 28749 17796
rect 34669 17796 34709 22073
rect 35080 22073 41080 22113
rect 35080 17796 35120 22073
rect 34669 16153 35120 17796
rect 41040 17796 41080 22073
rect 41451 22073 47451 22113
rect 41451 17796 41491 22073
rect 41040 16153 41491 17796
rect 47411 17796 47451 22073
rect 47822 22073 53822 22113
rect 47822 17796 47862 22073
rect 47411 16153 47862 17796
rect 53782 17796 53822 22073
rect 54193 22073 60193 22113
rect 54193 17796 54233 22073
rect 53782 16153 54233 17796
rect 60153 17796 60193 22073
rect 60153 16153 60524 17796
rect -3186 16113 60524 16153
rect -3146 15742 -1463 16113
rect 3225 15742 4908 16113
rect 9596 15742 11279 16113
rect 15967 15742 17650 16113
rect 22338 15742 24021 16113
rect 28709 15742 30392 16113
rect 35080 15742 36763 16113
rect 41451 15742 43134 16113
rect 47822 15742 49505 16113
rect 54193 15742 55876 16113
rect -3146 15702 2854 15742
rect -3146 11425 -3106 15702
rect -3186 9782 -3106 11425
rect 2814 11425 2854 15702
rect 3225 15702 9225 15742
rect 3225 11425 3265 15702
rect 2814 9782 3265 11425
rect 9185 11425 9225 15702
rect 9596 15702 15596 15742
rect 9596 11425 9636 15702
rect 9185 9782 9636 11425
rect 15556 11425 15596 15702
rect 15967 15702 21967 15742
rect 15967 11425 16007 15702
rect 15556 9782 16007 11425
rect 21927 11425 21967 15702
rect 22338 15702 28338 15742
rect 22338 11425 22378 15702
rect 21927 9782 22378 11425
rect 28298 11425 28338 15702
rect 28709 15702 34709 15742
rect 28709 11425 28749 15702
rect 28298 9782 28749 11425
rect 34669 11425 34709 15702
rect 35080 15702 41080 15742
rect 35080 11425 35120 15702
rect 34669 9782 35120 11425
rect 41040 11425 41080 15702
rect 41451 15702 47451 15742
rect 41451 11425 41491 15702
rect 41040 9782 41491 11425
rect 47411 11425 47451 15702
rect 47822 15702 53822 15742
rect 47822 11425 47862 15702
rect 47411 9782 47862 11425
rect 53782 11425 53822 15702
rect 54193 15702 60193 15742
rect 54193 11425 54233 15702
rect 53782 9782 54233 11425
rect 60153 11425 60193 15702
rect 60153 9782 60524 11425
rect -3186 9742 60524 9782
rect -3146 9371 -1463 9742
rect 3225 9371 4908 9742
rect 9596 9371 11279 9742
rect 15967 9371 17650 9742
rect 22338 9371 24021 9742
rect 28709 9371 30392 9742
rect 35080 9371 36763 9742
rect 41451 9371 43134 9742
rect 47822 9371 49505 9742
rect 54193 9371 55876 9742
rect -3146 9331 2854 9371
rect -3146 5054 -3106 9331
rect -3186 3411 -3106 5054
rect 2814 5054 2854 9331
rect 3225 9331 9225 9371
rect 3225 5054 3265 9331
rect 2814 3411 3265 5054
rect 9185 5054 9225 9331
rect 9596 9331 15596 9371
rect 9596 5054 9636 9331
rect 9185 3411 9636 5054
rect 15556 5054 15596 9331
rect 15967 9331 21967 9371
rect 15967 5054 16007 9331
rect 15556 3411 16007 5054
rect 21927 5054 21967 9331
rect 22338 9331 28338 9371
rect 22338 5054 22378 9331
rect 21927 3411 22378 5054
rect 28298 5054 28338 9331
rect 28709 9331 34709 9371
rect 28709 5054 28749 9331
rect 28298 3411 28749 5054
rect 34669 5054 34709 9331
rect 35080 9331 41080 9371
rect 35080 5054 35120 9331
rect 34669 3411 35120 5054
rect 41040 5054 41080 9331
rect 41451 9331 47451 9371
rect 41451 5054 41491 9331
rect 41040 3411 41491 5054
rect 47411 5054 47451 9331
rect 47822 9331 53822 9371
rect 47822 5054 47862 9331
rect 47411 3411 47862 5054
rect 53782 5054 53822 9331
rect 54193 9331 60193 9371
rect 54193 5054 54233 9331
rect 53782 3411 54233 5054
rect 60153 5054 60193 9331
rect 60153 3411 60524 5054
rect -3186 3371 60524 3411
rect -3146 3000 -1463 3371
rect 3225 3000 4908 3371
rect 9596 3000 11279 3371
rect 15967 3000 17650 3371
rect 22338 3000 24021 3371
rect 28709 3000 30392 3371
rect 35080 3000 36763 3371
rect 41451 3000 43134 3371
rect 47822 3000 49505 3371
rect 54193 3000 55876 3371
rect -3146 2960 2854 3000
rect -3146 -1317 -3106 2960
rect -3186 -2960 -3106 -1317
rect 2814 -1317 2854 2960
rect 3225 2960 9225 3000
rect 3225 -1317 3265 2960
rect 2814 -2960 3265 -1317
rect 9185 -1317 9225 2960
rect 9596 2960 15596 3000
rect 9596 -1317 9636 2960
rect 9185 -2960 9636 -1317
rect 15556 -1317 15596 2960
rect 15967 2960 21967 3000
rect 15967 -1317 16007 2960
rect 15556 -2960 16007 -1317
rect 21927 -1317 21967 2960
rect 22338 2960 28338 3000
rect 22338 -1317 22378 2960
rect 21927 -2960 22378 -1317
rect 28298 -1317 28338 2960
rect 28709 2960 34709 3000
rect 28709 -1317 28749 2960
rect 28298 -2960 28749 -1317
rect 34669 -1317 34709 2960
rect 35080 2960 41080 3000
rect 35080 -1317 35120 2960
rect 34669 -2960 35120 -1317
rect 41040 -1317 41080 2960
rect 41451 2960 47451 3000
rect 41451 -1317 41491 2960
rect 41040 -2960 41491 -1317
rect 47411 -1317 47451 2960
rect 47822 2960 53822 3000
rect 47822 -1317 47862 2960
rect 47411 -2960 47862 -1317
rect 53782 -1317 53822 2960
rect 54193 2960 60193 3000
rect 54193 -1317 54233 2960
rect 53782 -2960 54233 -1317
rect 60153 -1317 60193 2960
rect 60153 -2960 60524 -1317
rect -3186 -3000 60524 -2960
rect -3146 -3040 -1463 -3000
rect 3225 -3040 4908 -3000
rect 9596 -3040 11279 -3000
rect 15967 -3040 17650 -3000
rect 22338 -3040 24021 -3000
rect 28709 -3040 30392 -3000
rect 35080 -3040 36763 -3000
rect 41451 -3040 43134 -3000
rect 47822 -3040 49505 -3000
rect 54193 -3040 55876 -3000
<< properties >>
string FIXED_BBOX -3186 -3040 2894 3040
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 30 l 30 val 1.822k carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
