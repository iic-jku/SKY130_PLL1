magic
tech sky130A
magscale 1 2
timestamp 1666529776
<< error_s >>
rect 2817 1245 2875 1251
rect 2817 1211 2829 1245
rect 2817 1205 2875 1211
rect 3246 992 3255 999
rect 3297 992 3306 999
rect 3246 990 3250 992
rect 3302 990 3306 992
rect 1185 977 1243 983
rect 3237 981 3246 990
rect 3306 981 3315 990
rect 1185 943 1197 977
rect 1185 937 1243 943
rect 3237 930 3246 939
rect 3306 930 3315 939
rect 3246 928 3250 930
rect 3302 928 3306 930
rect 3246 921 3255 928
rect 3297 921 3306 928
<< locali >>
rect 1277 1205 2015 1251
rect 2429 1205 2591 1251
rect 2045 937 2399 983
rect 2621 937 2783 983
<< metal1 >>
rect 2056 2309 2126 2315
rect 2056 1717 2126 2239
rect -154 1647 929 1717
rect 999 1647 3869 1717
rect 3939 1647 3945 1717
rect 1949 1553 2019 1559
rect -154 1483 -27 1553
rect 43 1483 1949 1553
rect 2019 1483 2915 1553
rect 2985 1483 2991 1553
rect 3061 1453 3131 1647
rect 2484 1441 2536 1447
rect 2484 1383 2536 1389
rect 462 1202 468 1254
rect 520 1251 526 1254
rect 2489 1251 2531 1383
rect 3061 1377 3131 1383
rect 520 1205 2015 1251
rect 2429 1205 2591 1251
rect 520 1202 526 1205
rect 3244 983 3250 986
rect 2045 937 2399 983
rect 2621 937 3250 983
rect 2201 826 2243 937
rect 3244 934 3250 937
rect 3302 934 3308 986
rect 3495 826 3501 831
rect 2201 784 3501 826
rect 3495 779 3501 784
rect 3553 779 3559 831
rect 1965 634 2337 668
rect 3056 253 3108 259
rect -95 206 -53 248
rect 2119 201 2125 253
rect 2177 201 2183 253
rect 3056 195 3108 201
rect 1773 -195 2433 -161
rect 3061 -375 3103 195
<< via1 >>
rect 2056 2239 2126 2309
rect 929 1647 999 1717
rect 3869 1647 3939 1717
rect -27 1483 43 1553
rect 1949 1483 2019 1553
rect 2915 1483 2985 1553
rect 2484 1389 2536 1441
rect 3061 1383 3131 1453
rect 468 1202 520 1254
rect 3250 934 3302 986
rect 3501 779 3553 831
rect 2125 201 2177 253
rect 3056 201 3108 253
<< metal2 >>
rect 464 3001 524 3010
rect 464 2932 524 2941
rect 3658 3001 3718 3010
rect 3658 2932 3718 2941
rect 473 2908 515 2932
rect 3667 2908 3709 2932
rect 1826 2619 2356 2689
rect 2056 2309 2126 2619
rect 2050 2239 2056 2309
rect 2126 2239 2132 2309
rect 1730 1980 2452 2050
rect -27 1553 43 1559
rect -27 -53 43 1483
rect 473 1260 515 1812
rect 929 1717 999 1723
rect 468 1254 520 1260
rect 468 1196 520 1202
rect 929 1164 999 1647
rect 1949 1553 2019 1980
rect 3667 1703 3709 1812
rect 1949 1477 2019 1483
rect 2489 1661 3709 1703
rect 3869 1717 3939 1723
rect 2489 1441 2531 1661
rect 3939 1647 4425 1717
rect 3869 1641 3939 1647
rect 4355 1579 4425 1647
rect 2915 1553 2985 1559
rect 2985 1483 3786 1553
rect 2915 1477 2985 1483
rect 2478 1389 2484 1441
rect 2536 1389 2542 1441
rect 3055 1383 3061 1453
rect 3131 1383 3137 1453
rect 3061 1164 3131 1383
rect 929 1094 1137 1164
rect 2923 1094 3131 1164
rect 929 586 999 1094
rect 2475 585 2545 996
rect 3250 990 3302 992
rect 3250 928 3302 930
rect 2125 253 2177 259
rect 3050 201 3056 253
rect 3108 201 3114 253
rect 2125 195 2177 201
rect 3398 -53 3468 1483
rect 3501 831 3553 837
rect 3501 773 3553 779
rect 3506 226 3548 773
rect 4677 277 4737 286
rect 4644 226 4677 268
rect 4677 208 4737 217
rect -27 -123 181 -53
rect 1822 -123 2385 -53
rect 2827 -123 3468 -53
<< via2 >>
rect 464 2941 524 3001
rect 3658 2941 3718 3001
rect 3246 986 3306 990
rect 3246 934 3250 986
rect 3250 934 3302 986
rect 3302 934 3306 986
rect 3246 930 3306 934
rect 4677 217 4737 277
<< metal3 >>
rect 459 3001 529 3006
rect 3653 3001 3723 3006
rect 459 2941 464 3001
rect 524 2941 3658 3001
rect 3718 2941 4737 3001
rect 459 2936 529 2941
rect 3653 2936 3723 2941
rect 3241 990 3311 995
rect 4677 990 4737 2941
rect 3241 930 3246 990
rect 3306 930 4737 990
rect 3241 925 3311 930
rect 4677 282 4737 930
rect 4672 277 4742 282
rect 4672 217 4677 277
rect 4737 217 4742 277
rect 4672 212 4742 217
use buffer  buffer_0
timestamp 1666523630
transform 1 0 -53 0 1 -333
box 0 0 2204 1138
use simple_inv  simple_inv_0
timestamp 1666523630
transform 1 0 2204 0 1 280
box -53 -613 857 525
use cap50f  sky130_fd_pr__cap_mim_m3_1_H9XL9H_0
timestamp 1666529717
transform 1 0 2511 0 1 -933
box -650 -600 649 600
use slope_p  sky130_fd_pr__pfet_01v8_BDAFKN_0
timestamp 1666523630
transform 1 0 2030 0 1 1094
box -1031 -289 1031 289
use tgate_1  tgate_1_0
timestamp 1666523630
transform 0 -1 1054 -1 0 2689
box -261 -952 919 1138
use tgate_1  tgate_1_1
timestamp 1666523630
transform 0 1 3128 -1 0 2689
box -261 -952 919 1138
use tgate_1  tgate_1_2
timestamp 1666523630
transform -1 0 4425 0 -1 807
box -261 -952 919 1138
<< labels >>
rlabel metal1 -95 206 -53 248 0 clk_in
rlabel metal1 3061 -375 3103 -333 5 clk_out
rlabel metal3 4677 930 4737 990 0 v_bias
rlabel metal1 -154 1647 -84 1717 3 vdd
rlabel metal1 -154 1483 -84 1553 0 vss
rlabel space 1964 2908 2006 2950 0 bit2
rlabel space 2176 2908 2218 2950 3 bit0
rlabel space 4644 1717 4686 1759 0 bit1
<< end >>
