magic
tech sky130A
magscale 1 2
timestamp 1668357910
<< pwell >>
rect -359 -280 359 280
<< nmos >>
rect -159 -70 -129 70
rect -63 -70 -33 70
rect 33 -70 63 70
rect 129 -70 159 70
<< ndiff >>
rect -221 58 -159 70
rect -221 -58 -209 58
rect -175 -58 -159 58
rect -221 -70 -159 -58
rect -129 58 -63 70
rect -129 -58 -113 58
rect -79 -58 -63 58
rect -129 -70 -63 -58
rect -33 58 33 70
rect -33 -58 -17 58
rect 17 -58 33 58
rect -33 -70 33 -58
rect 63 58 129 70
rect 63 -58 79 58
rect 113 -58 129 58
rect 63 -70 129 -58
rect 159 58 221 70
rect 159 -58 175 58
rect 209 -58 221 58
rect 159 -70 221 -58
<< ndiffc >>
rect -209 -58 -175 58
rect -113 -58 -79 58
rect -17 -58 17 58
rect 79 -58 113 58
rect 175 -58 209 58
<< psubdiff >>
rect -323 210 -227 244
rect 227 210 323 244
rect -323 148 -289 210
rect 289 148 323 210
rect -323 -210 -289 -148
rect 289 -210 323 -148
rect -323 -244 -227 -210
rect 227 -244 323 -210
<< psubdiffcont >>
rect -227 210 227 244
rect -323 -148 -289 148
rect 289 -148 323 148
rect -227 -244 227 -210
<< poly >>
rect -177 142 -111 158
rect -177 108 -161 142
rect -127 108 -111 142
rect -177 92 -111 108
rect 111 142 177 158
rect 111 108 127 142
rect 161 108 177 142
rect -159 70 -129 92
rect -63 70 -33 96
rect 33 70 63 96
rect 111 92 177 108
rect 129 70 159 92
rect -159 -96 -129 -70
rect -63 -92 -33 -70
rect 33 -92 63 -70
rect -81 -108 81 -92
rect 129 -96 159 -70
rect -81 -142 -65 -108
rect -31 -142 31 -108
rect 65 -142 81 -108
rect -81 -158 81 -142
<< polycont >>
rect -161 108 -127 142
rect 127 108 161 142
rect -65 -142 -31 -108
rect 31 -142 65 -108
<< locali >>
rect -323 210 -227 244
rect 227 210 323 244
rect -323 148 -289 210
rect 289 148 323 210
rect -177 108 -161 142
rect -127 108 -111 142
rect 111 108 127 142
rect 161 108 177 142
rect -209 58 -175 74
rect -209 -74 -175 -58
rect -113 58 -79 74
rect -113 -74 -79 -58
rect -17 58 17 74
rect -17 -74 17 -58
rect 79 58 113 74
rect 79 -74 113 -58
rect 175 58 209 74
rect 175 -74 209 -58
rect -81 -142 -65 -108
rect -31 -142 31 -108
rect 65 -142 81 -108
rect -323 -210 -289 -148
rect 289 -210 323 -148
rect -323 -244 -227 -210
rect 227 -244 323 -210
<< viali >>
rect -161 108 -127 142
rect 127 108 161 142
rect -209 -58 -175 58
rect -113 -58 -79 58
rect -17 -58 17 58
rect 79 -58 113 58
rect 175 -58 209 58
rect -65 -142 -31 -108
rect 31 -142 65 -108
<< metal1 >>
rect -209 142 -115 148
rect -209 108 -161 142
rect -127 108 -115 142
rect -209 102 -115 108
rect 115 142 209 148
rect 115 108 127 142
rect 161 108 209 142
rect 115 102 209 108
rect -209 70 -173 102
rect 173 70 209 102
rect -215 58 -169 70
rect -215 0 -209 58
rect -220 -7 -209 0
rect -175 0 -169 58
rect -119 58 -73 70
rect -119 0 -113 58
rect -175 -7 -113 0
rect -79 0 -73 58
rect -23 58 23 70
rect -79 -7 -68 0
rect -220 -63 -218 -7
rect -165 -63 -122 -7
rect -69 -63 -68 -7
rect -220 -70 -68 -63
rect -23 -58 -17 58
rect 17 -58 23 58
rect 73 58 119 70
rect 73 0 79 58
rect -23 -70 23 -58
rect 68 -7 79 0
rect 113 0 119 58
rect 169 58 215 70
rect 169 0 175 58
rect 113 -7 175 0
rect 209 0 215 58
rect 209 -7 220 0
rect 68 -63 69 -7
rect 122 -63 165 -7
rect 218 -63 220 -7
rect 68 -70 220 -63
rect -77 -108 77 -102
rect -77 -142 -65 -108
rect -31 -142 31 -108
rect 65 -142 77 -108
rect -77 -148 77 -142
<< via1 >>
rect -218 -58 -209 -7
rect -209 -58 -175 -7
rect -175 -58 -165 -7
rect -218 -63 -165 -58
rect -122 -58 -113 -7
rect -113 -58 -79 -7
rect -79 -58 -69 -7
rect -122 -63 -69 -58
rect 69 -58 79 -7
rect 79 -58 113 -7
rect 113 -58 122 -7
rect 69 -63 122 -58
rect 165 -58 175 -7
rect 175 -58 209 -7
rect 209 -58 218 -7
rect 165 -63 218 -58
<< metal2 >>
rect -220 -7 -68 0
rect -220 -63 -218 -7
rect -165 -63 -122 -7
rect -69 -28 -68 -7
rect 68 -7 220 0
rect 68 -28 69 -7
rect -69 -63 69 -28
rect 122 -63 165 -7
rect 218 -63 220 -7
rect -220 -70 220 -63
<< properties >>
string FIXED_BBOX -306 -227 306 227
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.7 l 0.150 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
