magic
tech sky130A
magscale 1 2
timestamp 1668438816
<< locali >>
rect 628 2666 787 3063
<< viali >>
rect 787 2666 1184 3063
<< metal1 >>
rect 112 3063 512 3080
rect 112 2666 129 3063
rect 497 2666 512 3063
rect 112 2650 512 2666
rect 781 3069 1190 3075
rect 781 3063 793 3069
rect 781 2666 787 3063
rect 781 2660 793 2666
rect 1190 2660 1196 3069
rect 781 2654 1190 2660
rect 114 528 514 544
rect 114 130 128 528
rect 498 130 514 528
rect 114 112 514 130
<< via1 >>
rect 129 2666 497 3063
rect 793 3063 1190 3069
rect 793 2666 1184 3063
rect 1184 2666 1190 3063
rect 793 2660 1190 2666
rect 128 130 498 528
<< metal2 >>
rect 112 3063 512 3080
rect 793 3069 1190 3075
rect 112 2666 129 3063
rect 497 2666 512 3063
rect 112 2650 512 2666
rect 784 2660 793 3069
rect 1190 2660 1199 3069
rect 793 2654 1190 2660
rect 114 528 514 544
rect 114 130 128 528
rect 498 130 514 528
rect 114 112 514 130
<< via2 >>
rect 793 2660 1190 3069
<< metal3 >>
rect 788 3069 798 3074
rect 788 2660 793 3069
rect 788 2655 798 2660
rect 1195 2655 1201 3074
<< via3 >>
rect 798 3069 1195 3074
rect 798 2660 1190 3069
rect 1190 2660 1195 3069
rect 798 2655 1195 2660
<< metal4 >>
rect 797 3074 799 3075
rect 797 2655 798 3074
rect 797 2654 799 2655
<< via4 >>
rect 799 3074 1196 3075
rect 799 2655 1195 3074
rect 1195 2655 1196 3074
rect 799 2654 1196 2655
<< metal5 >>
rect 775 3075 1220 3099
rect 775 2654 799 3075
rect 1196 2654 1220 3075
rect 775 2630 1220 2654
use sky130_fd_pr__res_generic_po_PL36XQ  sky130_fd_pr__res_generic_po_PL36XQ_0
timestamp 1668438816
transform 1 0 313 0 1 1596
box -366 -1649 366 1649
<< end >>
