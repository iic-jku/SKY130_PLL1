magic
tech sky130A
magscale 1 2
timestamp 1668153059
<< xpolycontact >>
rect 113 4881 683 5313
rect 13201 4881 13771 5313
rect 5021 4117 5591 4549
rect 6657 4117 7227 4549
rect 8293 4117 8863 4549
rect 9929 4117 10499 4549
rect 11565 4117 12135 4549
rect 13201 4117 13771 4549
<< metal1 >>
rect 12383 9287 12953 10023
rect 931 9269 1501 9287
rect 931 8872 947 9269
rect 1485 8872 1501 9269
rect 931 8855 1501 8872
rect 1749 9269 3137 9287
rect 1749 8872 2583 9269
rect 3121 8872 3137 9269
rect 1749 8855 3137 8872
rect 3385 9269 4773 9287
rect 3385 8872 4219 9269
rect 4757 8872 4773 9269
rect 3385 8855 4773 8872
rect 5021 9269 6409 9287
rect 5021 8872 5855 9269
rect 6393 8872 6409 9269
rect 5021 8855 6409 8872
rect 6657 9269 8045 9287
rect 6657 8872 7491 9269
rect 8029 8872 8045 9269
rect 6657 8855 8045 8872
rect 8293 9269 9681 9287
rect 8293 8872 9127 9269
rect 9665 8872 9681 9269
rect 8293 8855 9681 8872
rect 9929 9269 11317 9287
rect 9929 8872 10763 9269
rect 11301 8872 11317 9269
rect 9929 8855 11317 8872
rect 11565 8855 12953 9287
rect 113 5295 683 5313
rect 113 4898 129 5295
rect 667 4898 683 5295
rect 113 4881 683 4898
rect 931 4117 1501 5313
rect 1749 5296 2319 5313
rect 1749 4899 1765 5296
rect 2303 4899 2319 5296
rect 1749 4117 2319 4899
rect 2567 4117 3137 5313
rect 3385 4531 3955 4549
rect 3385 4134 3401 4531
rect 3939 4134 3955 4531
rect 3385 4117 3955 4134
rect 4203 4117 4773 5313
rect 5021 4531 5591 4549
rect 5021 4134 5037 4531
rect 5575 4134 5591 4531
rect 5021 4117 5591 4134
rect 5839 4117 6409 5313
rect 6657 4531 7227 4549
rect 6657 4134 6673 4531
rect 7211 4134 7227 4531
rect 6657 4117 7227 4134
rect 7475 4117 8045 5313
rect 8293 4531 8863 4549
rect 8293 4134 8309 4531
rect 8847 4134 8863 4531
rect 8293 4117 8863 4134
rect 9111 4117 9681 5313
rect 9929 4531 10499 4549
rect 9929 4134 9945 4531
rect 10483 4134 10499 4531
rect 9929 4117 10499 4134
rect 10747 4117 11317 5313
rect 11565 4531 12135 4549
rect 11565 4134 11581 4531
rect 12119 4134 12135 4531
rect 11565 4117 12135 4134
rect 12383 4117 12953 5313
rect 13201 5295 13771 5313
rect 13201 4898 13217 5295
rect 13755 4898 13771 5295
rect 13201 4881 13771 4898
rect 13201 4531 13771 4549
rect 13201 4134 13217 4531
rect 13755 4134 13771 4531
rect 13201 4117 13771 4134
rect 1749 558 2319 575
rect 931 -593 1501 167
rect 1749 161 1765 558
rect 2303 161 2319 558
rect 3385 558 3955 575
rect 1749 143 2319 161
rect 2567 -593 3137 179
rect 3385 161 3401 558
rect 3939 161 3955 558
rect 3385 143 3955 161
rect 4203 -593 4773 167
rect 5839 -593 6409 176
rect 7475 -593 8045 176
rect 9111 -593 9681 175
rect 10747 -593 11317 175
rect 12383 -593 12953 175
<< via1 >>
rect 947 8872 1485 9269
rect 2583 8872 3121 9269
rect 4219 8872 4757 9269
rect 5855 8872 6393 9269
rect 7491 8872 8029 9269
rect 9127 8872 9665 9269
rect 10763 8872 11301 9269
rect 129 4898 667 5295
rect 1765 4899 2303 5296
rect 3401 4899 3939 5296
rect 3401 4134 3939 4531
rect 5037 4899 5575 5296
rect 5037 4134 5575 4531
rect 6673 4899 7211 5296
rect 6673 4134 7211 4531
rect 8309 4899 8847 5296
rect 8309 4134 8847 4531
rect 9945 4899 10483 5296
rect 9945 4134 10483 4531
rect 11581 4899 12119 5296
rect 11581 4134 12119 4531
rect 13217 4898 13755 5295
rect 13217 4134 13755 4531
rect 1765 161 2303 558
rect 3401 161 3939 558
<< metal2 >>
rect 931 9269 1501 9287
rect 931 8872 947 9269
rect 1485 8872 1501 9269
rect 931 5313 1501 8872
rect 2567 9269 3137 9287
rect 2567 8872 2583 9269
rect 3121 8872 3137 9269
rect 2567 5313 3137 8872
rect 4203 9269 4773 9287
rect 4203 8872 4219 9269
rect 4757 8872 4773 9269
rect 4203 5313 4773 8872
rect 5839 9269 6409 9287
rect 5839 8872 5855 9269
rect 6393 8872 6409 9269
rect 5839 5313 6409 8872
rect 7475 9269 8045 9287
rect 7475 8872 7491 9269
rect 8029 8872 8045 9269
rect 7475 5313 8045 8872
rect 9111 9269 9681 9287
rect 9111 8872 9127 9269
rect 9665 8872 9681 9269
rect 9111 5313 9681 8872
rect 10747 9269 11317 9287
rect 10747 8872 10763 9269
rect 11301 8872 11317 9269
rect 10747 5313 11317 8872
rect 113 5295 683 5313
rect 113 4898 129 5295
rect 667 4898 683 5295
rect 113 4549 683 4898
rect 931 5296 2319 5313
rect 931 4899 1765 5296
rect 2303 4899 2319 5296
rect 931 4881 2319 4899
rect 2567 5296 3955 5313
rect 2567 4899 3401 5296
rect 3939 4899 3955 5296
rect 2567 4881 3955 4899
rect 4203 5296 5591 5313
rect 4203 4899 5037 5296
rect 5575 4899 5591 5296
rect 4203 4881 5591 4899
rect 5839 5296 7227 5313
rect 5839 4899 6673 5296
rect 7211 4899 7227 5296
rect 5839 4881 7227 4899
rect 7475 5296 8863 5313
rect 7475 4899 8309 5296
rect 8847 4899 8863 5296
rect 7475 4881 8863 4899
rect 9111 5296 10499 5313
rect 9111 4899 9945 5296
rect 10483 4899 10499 5296
rect 9111 4881 10499 4899
rect 10747 5296 12135 5313
rect 10747 4899 11581 5296
rect 12119 4899 12135 5296
rect 10747 4881 12135 4899
rect 13201 5295 13771 5313
rect 13201 4898 13217 5295
rect 13755 4898 13771 5295
rect 13201 4549 13771 4898
rect -485 4531 13771 4549
rect -485 4134 3401 4531
rect 3939 4134 5037 4531
rect 5575 4134 6673 4531
rect 7211 4134 8309 4531
rect 8847 4134 9945 4531
rect 10483 4134 11581 4531
rect 12119 4134 13217 4531
rect 13755 4134 13771 4531
rect -485 4117 13771 4134
rect 1749 558 3955 575
rect 1749 161 1765 558
rect 2303 161 3401 558
rect 3939 161 3955 558
rect 1749 143 3955 161
use sky130_fd_pr__res_high_po_2p85_DZGNGK  sky130_fd_pr__res_high_po_2p85_DZGNGK_0
timestamp 1668153059
transform 1 0 6942 0 1 2346
box -6995 -2369 6995 2369
use sky130_fd_pr__res_high_po_2p85_DZGNGK  sky130_fd_pr__res_high_po_2p85_DZGNGK_1
timestamp 1668153059
transform 1 0 6942 0 1 7084
box -6995 -2369 6995 2369
<< labels >>
rlabel metal1 12383 9453 12953 10023 0 vout
rlabel metal1 931 -593 1501 -23 3 b0
rlabel metal1 2567 -593 3137 -23 3 b1
rlabel metal1 4203 -593 4773 -23 0 b2
rlabel metal1 5839 -593 6409 -23 5 b3
rlabel metal1 7475 -593 8045 -23 0 b4
rlabel metal1 9111 -593 9681 -23 0 b5
rlabel metal1 10747 -593 11317 -23 0 b6
rlabel metal1 12383 -593 12953 -23 0 b7
rlabel metal2 -485 4117 -53 4549 7 vss
<< end >>
