magic
tech sky130A
magscale 1 2
timestamp 1663426905
<< error_p >>
rect -653 151 -595 157
rect 595 151 653 157
rect -653 117 -641 151
rect 595 117 607 151
rect -653 111 -595 117
rect 595 111 653 117
<< nwell >>
rect -839 -289 839 289
<< pmos >>
rect -639 -70 -609 70
rect -543 -70 -513 70
rect -447 -70 -417 70
rect -351 -70 -321 70
rect -255 -70 -225 70
rect -159 -70 -129 70
rect -63 -70 -33 70
rect 33 -70 63 70
rect 129 -70 159 70
rect 225 -70 255 70
rect 321 -70 351 70
rect 417 -70 447 70
rect 513 -70 543 70
rect 609 -70 639 70
<< pdiff >>
rect -701 58 -639 70
rect -701 -58 -689 58
rect -655 -58 -639 58
rect -701 -70 -639 -58
rect -609 58 -543 70
rect -609 -58 -593 58
rect -559 -58 -543 58
rect -609 -70 -543 -58
rect -513 58 -447 70
rect -513 -58 -497 58
rect -463 -58 -447 58
rect -513 -70 -447 -58
rect -417 58 -351 70
rect -417 -58 -401 58
rect -367 -58 -351 58
rect -417 -70 -351 -58
rect -321 58 -255 70
rect -321 -58 -305 58
rect -271 -58 -255 58
rect -321 -70 -255 -58
rect -225 58 -159 70
rect -225 -58 -209 58
rect -175 -58 -159 58
rect -225 -70 -159 -58
rect -129 58 -63 70
rect -129 -58 -113 58
rect -79 -58 -63 58
rect -129 -70 -63 -58
rect -33 58 33 70
rect -33 -58 -17 58
rect 17 -58 33 58
rect -33 -70 33 -58
rect 63 58 129 70
rect 63 -58 79 58
rect 113 -58 129 58
rect 63 -70 129 -58
rect 159 58 225 70
rect 159 -58 175 58
rect 209 -58 225 58
rect 159 -70 225 -58
rect 255 58 321 70
rect 255 -58 271 58
rect 305 -58 321 58
rect 255 -70 321 -58
rect 351 58 417 70
rect 351 -58 367 58
rect 401 -58 417 58
rect 351 -70 417 -58
rect 447 58 513 70
rect 447 -58 463 58
rect 497 -58 513 58
rect 447 -70 513 -58
rect 543 58 609 70
rect 543 -58 559 58
rect 593 -58 609 58
rect 543 -70 609 -58
rect 639 58 701 70
rect 639 -58 655 58
rect 689 -58 701 58
rect 639 -70 701 -58
<< pdiffc >>
rect -689 -58 -655 58
rect -593 -58 -559 58
rect -497 -58 -463 58
rect -401 -58 -367 58
rect -305 -58 -271 58
rect -209 -58 -175 58
rect -113 -58 -79 58
rect -17 -58 17 58
rect 79 -58 113 58
rect 175 -58 209 58
rect 271 -58 305 58
rect 367 -58 401 58
rect 463 -58 497 58
rect 559 -58 593 58
rect 655 -58 689 58
<< nsubdiff >>
rect -803 219 -707 253
rect 707 219 803 253
rect -803 157 -769 219
rect 769 157 803 219
rect -803 -219 -769 -157
rect 769 -219 803 -157
rect -803 -253 -707 -219
rect 707 -253 803 -219
<< nsubdiffcont >>
rect -707 219 707 253
rect -803 -157 -769 157
rect 769 -157 803 157
rect -707 -253 707 -219
<< poly >>
rect -657 151 -591 167
rect -657 117 -641 151
rect -607 117 -591 151
rect -657 101 -591 117
rect 591 151 657 167
rect 591 117 607 151
rect 641 117 657 151
rect 591 101 657 117
rect -639 70 -609 101
rect -543 70 -513 96
rect -447 70 -417 96
rect -351 70 -321 96
rect -255 70 -225 96
rect -159 70 -129 96
rect -63 70 -33 96
rect 33 70 63 96
rect 129 70 159 96
rect 225 70 255 96
rect 321 70 351 96
rect 417 70 447 96
rect 513 70 543 96
rect 609 70 639 101
rect -639 -96 -609 -70
rect -543 -101 -513 -70
rect -447 -101 -417 -70
rect -351 -101 -321 -70
rect -255 -101 -225 -70
rect -159 -101 -129 -70
rect -63 -101 -33 -70
rect 33 -101 63 -70
rect 129 -101 159 -70
rect 225 -101 255 -70
rect 321 -101 351 -70
rect 417 -101 447 -70
rect 513 -101 543 -70
rect 609 -96 639 -70
rect -561 -117 561 -101
rect -561 -151 -545 -117
rect -511 -151 -449 -117
rect -415 -151 -353 -117
rect -319 -151 -257 -117
rect -223 -151 -161 -117
rect -127 -151 -65 -117
rect -31 -151 31 -117
rect 65 -151 127 -117
rect 161 -151 223 -117
rect 257 -151 319 -117
rect 353 -151 415 -117
rect 449 -151 511 -117
rect 545 -151 561 -117
rect -561 -167 561 -151
<< polycont >>
rect -641 117 -607 151
rect 607 117 641 151
rect -545 -151 -511 -117
rect -449 -151 -415 -117
rect -353 -151 -319 -117
rect -257 -151 -223 -117
rect -161 -151 -127 -117
rect -65 -151 -31 -117
rect 31 -151 65 -117
rect 127 -151 161 -117
rect 223 -151 257 -117
rect 319 -151 353 -117
rect 415 -151 449 -117
rect 511 -151 545 -117
<< locali >>
rect -803 219 -707 253
rect 707 219 803 253
rect -803 157 -769 219
rect 769 157 803 219
rect -657 117 -641 151
rect -607 117 -591 151
rect 591 117 607 151
rect 641 117 657 151
rect -689 58 -655 74
rect -689 -74 -655 -58
rect -593 58 -559 74
rect -593 -74 -559 -58
rect -497 58 -463 74
rect -497 -74 -463 -58
rect -401 58 -367 74
rect -401 -74 -367 -58
rect -305 58 -271 74
rect -305 -74 -271 -58
rect -209 58 -175 74
rect -209 -74 -175 -58
rect -113 58 -79 74
rect -113 -74 -79 -58
rect -17 58 17 74
rect -17 -74 17 -58
rect 79 58 113 74
rect 79 -74 113 -58
rect 175 58 209 74
rect 175 -74 209 -58
rect 271 58 305 74
rect 271 -74 305 -58
rect 367 58 401 74
rect 367 -74 401 -58
rect 463 58 497 74
rect 463 -74 497 -58
rect 559 58 593 74
rect 559 -74 593 -58
rect 655 58 689 74
rect 655 -74 689 -58
rect -561 -151 -545 -117
rect -511 -151 -449 -117
rect -415 -151 -353 -117
rect -319 -151 -257 -117
rect -223 -151 -161 -117
rect -127 -151 -65 -117
rect -31 -151 31 -117
rect 65 -151 127 -117
rect 161 -151 223 -117
rect 257 -151 319 -117
rect 353 -151 415 -117
rect 449 -151 511 -117
rect 545 -151 561 -117
rect -803 -219 -769 -157
rect 769 -219 803 -157
rect -803 -253 -707 -219
rect 707 -253 803 -219
<< viali >>
rect -641 117 -607 151
rect 607 117 641 151
rect -689 -58 -655 58
rect -593 -58 -559 58
rect -497 -58 -463 58
rect -401 -58 -367 58
rect -305 -58 -271 58
rect -209 -58 -175 58
rect -113 -58 -79 58
rect -17 -58 17 58
rect 79 -58 113 58
rect 175 -58 209 58
rect 271 -58 305 58
rect 367 -58 401 58
rect 463 -58 497 58
rect 559 -58 593 58
rect 655 -58 689 58
rect -545 -151 -511 -117
rect -449 -151 -415 -117
rect -353 -151 -319 -117
rect -257 -151 -223 -117
rect -161 -151 -127 -117
rect -65 -151 -31 -117
rect 31 -151 65 -117
rect 127 -151 161 -117
rect 223 -151 257 -117
rect 319 -151 353 -117
rect 415 -151 449 -117
rect 511 -151 545 -117
<< metal1 >>
rect -653 151 -595 157
rect -653 117 -641 151
rect -607 117 -595 151
rect -653 111 -595 117
rect 595 151 653 157
rect 595 117 607 151
rect 641 117 653 151
rect 595 111 653 117
rect -703 61 -641 70
rect -703 9 -698 61
rect -646 9 -641 61
rect -703 0 -689 9
rect -695 -58 -689 0
rect -655 0 -641 9
rect -607 61 -545 70
rect -607 9 -602 61
rect -550 9 -545 61
rect -607 0 -593 9
rect -655 -58 -649 0
rect -695 -70 -649 -58
rect -599 -58 -593 0
rect -559 0 -545 9
rect -503 58 -457 70
rect -503 0 -497 58
rect -559 -58 -553 0
rect -599 -70 -553 -58
rect -511 -9 -497 0
rect -463 0 -457 58
rect -415 61 -353 70
rect -415 9 -410 61
rect -358 9 -353 61
rect -415 0 -401 9
rect -463 -9 -449 0
rect -511 -61 -506 -9
rect -454 -61 -449 -9
rect -511 -70 -449 -61
rect -407 -58 -401 0
rect -367 0 -353 9
rect -311 58 -265 70
rect -311 0 -305 58
rect -367 -58 -361 0
rect -407 -70 -361 -58
rect -319 -9 -305 0
rect -271 0 -265 58
rect -223 61 -161 70
rect -223 9 -218 61
rect -166 9 -161 61
rect -223 0 -209 9
rect -271 -9 -257 0
rect -319 -61 -314 -9
rect -262 -61 -257 -9
rect -319 -70 -257 -61
rect -215 -58 -209 0
rect -175 0 -161 9
rect -119 58 -73 70
rect -119 0 -113 58
rect -175 -58 -169 0
rect -215 -70 -169 -58
rect -127 -9 -113 0
rect -79 0 -73 58
rect -31 61 31 70
rect -31 9 -26 61
rect 26 9 31 61
rect -31 0 -17 9
rect -79 -9 -65 0
rect -127 -61 -122 -9
rect -70 -61 -65 -9
rect -127 -70 -65 -61
rect -23 -58 -17 0
rect 17 0 31 9
rect 73 58 119 70
rect 73 0 79 58
rect 17 -58 23 0
rect -23 -70 23 -58
rect 65 -9 79 0
rect 113 0 119 58
rect 161 61 223 70
rect 161 9 166 61
rect 218 9 223 61
rect 161 0 175 9
rect 113 -9 127 0
rect 65 -61 70 -9
rect 122 -61 127 -9
rect 65 -70 127 -61
rect 169 -58 175 0
rect 209 0 223 9
rect 265 58 311 70
rect 265 0 271 58
rect 209 -58 215 0
rect 169 -70 215 -58
rect 257 -9 271 0
rect 305 0 311 58
rect 353 61 415 70
rect 353 9 358 61
rect 410 9 415 61
rect 353 0 367 9
rect 305 -9 319 0
rect 257 -61 262 -9
rect 314 -61 319 -9
rect 257 -70 319 -61
rect 361 -58 367 0
rect 401 0 415 9
rect 457 58 503 70
rect 457 0 463 58
rect 401 -58 407 0
rect 361 -70 407 -58
rect 449 -9 463 0
rect 497 0 503 58
rect 545 61 607 70
rect 545 9 550 61
rect 602 9 607 61
rect 545 0 559 9
rect 497 -9 511 0
rect 449 -61 454 -9
rect 506 -61 511 -9
rect 449 -70 511 -61
rect 553 -58 559 0
rect 593 0 607 9
rect 641 61 701 70
rect 641 9 646 61
rect 698 9 701 61
rect 641 0 655 9
rect 593 -58 599 0
rect 553 -70 599 -58
rect 649 -58 655 0
rect 689 0 701 9
rect 689 -58 695 0
rect 649 -70 695 -58
rect -557 -117 -499 -111
rect -461 -117 -403 -111
rect -365 -117 -307 -111
rect -269 -117 -211 -111
rect -173 -117 -115 -111
rect -77 -117 -19 -111
rect 19 -117 77 -111
rect 115 -117 173 -111
rect 211 -117 269 -111
rect 307 -117 365 -111
rect 403 -117 461 -111
rect 499 -117 557 -111
rect -557 -151 -545 -117
rect -511 -151 -449 -117
rect -415 -151 -353 -117
rect -319 -151 -257 -117
rect -223 -151 -161 -117
rect -127 -151 -65 -117
rect -31 -151 31 -117
rect 65 -151 127 -117
rect 161 -151 223 -117
rect 257 -151 319 -117
rect 353 -151 415 -117
rect 449 -151 511 -117
rect 545 -151 557 -117
rect -557 -157 -499 -151
rect -461 -157 -403 -151
rect -365 -157 -307 -151
rect -269 -157 -211 -151
rect -173 -157 -115 -151
rect -77 -157 -19 -151
rect 19 -157 77 -151
rect 115 -157 173 -151
rect 211 -157 269 -151
rect 307 -157 365 -151
rect 403 -157 461 -151
rect 499 -157 557 -151
<< via1 >>
rect -698 58 -646 61
rect -698 9 -689 58
rect -689 9 -655 58
rect -655 9 -646 58
rect -602 58 -550 61
rect -602 9 -593 58
rect -593 9 -559 58
rect -559 9 -550 58
rect -410 58 -358 61
rect -410 9 -401 58
rect -401 9 -367 58
rect -367 9 -358 58
rect -506 -58 -497 -9
rect -497 -58 -463 -9
rect -463 -58 -454 -9
rect -506 -61 -454 -58
rect -218 58 -166 61
rect -218 9 -209 58
rect -209 9 -175 58
rect -175 9 -166 58
rect -314 -58 -305 -9
rect -305 -58 -271 -9
rect -271 -58 -262 -9
rect -314 -61 -262 -58
rect -26 58 26 61
rect -26 9 -17 58
rect -17 9 17 58
rect 17 9 26 58
rect -122 -58 -113 -9
rect -113 -58 -79 -9
rect -79 -58 -70 -9
rect -122 -61 -70 -58
rect 166 58 218 61
rect 166 9 175 58
rect 175 9 209 58
rect 209 9 218 58
rect 70 -58 79 -9
rect 79 -58 113 -9
rect 113 -58 122 -9
rect 70 -61 122 -58
rect 358 58 410 61
rect 358 9 367 58
rect 367 9 401 58
rect 401 9 410 58
rect 262 -58 271 -9
rect 271 -58 305 -9
rect 305 -58 314 -9
rect 262 -61 314 -58
rect 550 58 602 61
rect 550 9 559 58
rect 559 9 593 58
rect 593 9 602 58
rect 454 -58 463 -9
rect 463 -58 497 -9
rect 497 -58 506 -9
rect 454 -61 506 -58
rect 646 58 698 61
rect 646 9 655 58
rect 655 9 689 58
rect 689 9 698 58
<< metal2 >>
rect -709 63 -539 72
rect -709 7 -700 63
rect -644 7 -604 63
rect -548 7 -539 63
rect -709 -2 -539 7
rect -421 63 -347 72
rect -421 7 -412 63
rect -356 7 -347 63
rect -511 -9 -449 0
rect -421 -2 -347 7
rect -229 63 -155 72
rect -229 7 -220 63
rect -164 7 -155 63
rect -511 -61 -506 -9
rect -454 -36 -449 -9
rect -319 -9 -257 0
rect -229 -2 -155 7
rect -37 63 37 72
rect -37 7 -28 63
rect 28 7 37 63
rect -319 -36 -314 -9
rect -454 -61 -314 -36
rect -262 -36 -257 -9
rect -127 -9 -65 0
rect -37 -2 37 7
rect 155 63 229 72
rect 155 7 164 63
rect 220 7 229 63
rect -127 -36 -122 -9
rect -262 -61 -122 -36
rect -70 -36 -65 -9
rect 65 -9 127 0
rect 155 -2 229 7
rect 347 63 421 72
rect 347 7 356 63
rect 412 7 421 63
rect 65 -36 70 -9
rect -70 -61 70 -36
rect 122 -36 127 -9
rect 257 -9 319 0
rect 347 -2 421 7
rect 539 63 709 72
rect 539 7 548 63
rect 604 7 644 63
rect 700 7 709 63
rect 257 -36 262 -9
rect 122 -61 262 -36
rect 314 -36 319 -9
rect 449 -9 511 0
rect 539 -2 709 7
rect 449 -36 454 -9
rect 314 -61 454 -36
rect 506 -61 511 -9
rect -511 -70 511 -61
<< via2 >>
rect -700 61 -644 63
rect -700 9 -698 61
rect -698 9 -646 61
rect -646 9 -644 61
rect -700 7 -644 9
rect -604 61 -548 63
rect -604 9 -602 61
rect -602 9 -550 61
rect -550 9 -548 61
rect -604 7 -548 9
rect -412 61 -356 63
rect -412 9 -410 61
rect -410 9 -358 61
rect -358 9 -356 61
rect -412 7 -356 9
rect -220 61 -164 63
rect -220 9 -218 61
rect -218 9 -166 61
rect -166 9 -164 61
rect -220 7 -164 9
rect -28 61 28 63
rect -28 9 -26 61
rect -26 9 26 61
rect 26 9 28 61
rect -28 7 28 9
rect 164 61 220 63
rect 164 9 166 61
rect 166 9 218 61
rect 218 9 220 61
rect 164 7 220 9
rect 356 61 412 63
rect 356 9 358 61
rect 358 9 410 61
rect 410 9 412 61
rect 356 7 412 9
rect 548 61 604 63
rect 548 9 550 61
rect 550 9 602 61
rect 602 9 604 61
rect 548 7 604 9
rect 644 61 700 63
rect 644 9 646 61
rect 646 9 698 61
rect 698 9 700 61
rect 644 7 700 9
<< metal3 >>
rect -709 70 -539 72
rect -421 70 -347 72
rect -229 70 -155 72
rect -37 70 37 72
rect 155 70 229 72
rect 347 70 421 72
rect 539 70 709 72
rect -709 63 709 70
rect -709 7 -700 63
rect -644 7 -604 63
rect -548 10 -412 63
rect -548 7 -539 10
rect -709 -2 -539 7
rect -421 7 -412 10
rect -356 10 -220 63
rect -356 7 -347 10
rect -421 -2 -347 7
rect -229 7 -220 10
rect -164 10 -28 63
rect -164 7 -155 10
rect -229 -2 -155 7
rect -37 7 -28 10
rect 28 10 164 63
rect 28 7 37 10
rect -37 -2 37 7
rect 155 7 164 10
rect 220 10 356 63
rect 220 7 229 10
rect 155 -2 229 7
rect 347 7 356 10
rect 412 10 548 63
rect 412 7 421 10
rect 347 -2 421 7
rect 539 7 548 10
rect 604 7 644 63
rect 700 7 709 63
rect 539 -2 709 7
<< properties >>
string FIXED_BBOX -786 -236 786 236
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.7 l 0.15 m 1 nf 14 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
