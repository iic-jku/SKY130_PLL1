magic
tech sky130A
magscale 1 2
timestamp 1666523630
<< metal1 >>
rect 381 -32 423 79
rect -53 -74 423 -32
rect 381 -185 423 -74
<< metal2 >>
rect 381 -32 423 166
rect 381 -74 857 -32
rect 381 -263 423 -74
use sinv_n  sky130_fd_pr__nfet_01v8_2AA63J_0
timestamp 1666523630
transform 1 0 402 0 1 -333
box -359 -280 359 280
use sinv_p  sky130_fd_pr__pfet_01v8_X6FFBL_0
timestamp 1666523630
transform 1 0 402 0 1 236
box -455 -289 455 289
<< end >>
