magic
tech sky130A
magscale 1 2
timestamp 1660030277
<< pwell >>
rect -455 -280 455 280
<< nmos >>
rect -255 -70 -225 70
rect -159 -70 -129 70
rect -63 -70 -33 70
rect 33 -70 63 70
rect 129 -70 159 70
rect 225 -70 255 70
<< ndiff >>
rect -321 58 -255 70
rect -321 -58 -305 58
rect -271 -58 -255 58
rect -321 -70 -255 -58
rect -225 58 -159 70
rect -225 -58 -209 58
rect -175 -58 -159 58
rect -225 -70 -159 -58
rect -129 58 -63 70
rect -129 -58 -113 58
rect -79 -58 -63 58
rect -129 -70 -63 -58
rect -33 58 33 70
rect -33 -58 -17 58
rect 17 -58 33 58
rect -33 -70 33 -58
rect 63 58 129 70
rect 63 -58 79 58
rect 113 -58 129 58
rect 63 -70 129 -58
rect 159 58 225 70
rect 159 -58 175 58
rect 209 -58 225 58
rect 159 -70 225 -58
rect 255 58 321 70
rect 255 -58 271 58
rect 305 -58 321 58
rect 255 -70 321 -58
<< ndiffc >>
rect -305 -58 -271 58
rect -209 -58 -175 58
rect -113 -58 -79 58
rect -17 -58 17 58
rect 79 -58 113 58
rect 175 -58 209 58
rect 271 -58 305 58
<< psubdiff >>
rect -419 210 -323 244
rect 323 210 419 244
rect -419 148 -385 210
rect 385 148 419 210
rect -419 -210 -385 -148
rect 385 -210 419 -148
rect -419 -244 -323 -210
rect 323 -244 419 -210
<< psubdiffcont >>
rect -323 210 323 244
rect -419 -148 -385 148
rect 385 -148 419 148
rect -323 -244 323 -210
<< poly >>
rect -274 146 -208 162
rect -274 112 -258 146
rect -224 112 -208 146
rect -274 96 -208 112
rect 207 146 273 162
rect 207 112 223 146
rect 257 112 273 146
rect 207 96 273 112
rect -255 70 -225 96
rect -159 70 -129 96
rect -63 70 -33 96
rect 33 70 63 96
rect 129 70 159 96
rect 225 70 255 96
rect -255 -96 -225 -70
rect -159 -92 -129 -70
rect -177 -108 -111 -92
rect -63 -108 -33 -70
rect -177 -142 -161 -108
rect -127 -142 -33 -108
rect 33 -108 63 -70
rect 129 -92 159 -70
rect 111 -108 177 -92
rect 225 -96 255 -70
rect 33 -142 127 -108
rect 161 -142 177 -108
rect -177 -158 -111 -142
rect 111 -158 177 -142
<< polycont >>
rect -258 112 -224 146
rect 223 112 257 146
rect -161 -142 -127 -108
rect 127 -142 161 -108
<< locali >>
rect -419 210 -323 244
rect 323 210 419 244
rect -419 148 -385 210
rect 385 148 419 210
rect -274 112 -258 146
rect -224 112 -208 146
rect 207 112 223 146
rect 257 112 273 146
rect -305 58 -271 74
rect -305 -74 -271 -58
rect -209 58 -175 74
rect -209 -74 -175 -58
rect -113 58 -79 74
rect -113 -74 -79 -58
rect -17 58 17 74
rect -17 -74 17 -58
rect 79 58 113 74
rect 79 -74 113 -58
rect 175 58 209 74
rect 175 -74 209 -58
rect 271 58 305 74
rect 271 -74 305 -58
rect -177 -142 -161 -108
rect -127 -142 -111 -108
rect 111 -142 127 -108
rect 161 -142 177 -108
rect -419 -210 -385 -148
rect 385 -210 419 -148
rect -419 -244 -323 -210
rect 323 -244 419 -210
<< viali >>
rect -258 112 -224 146
rect 223 112 257 146
rect -305 -58 -271 58
rect -209 -58 -175 58
rect -113 -58 -79 58
rect -17 -58 17 58
rect 79 -58 113 58
rect 175 -58 209 58
rect 271 -58 305 58
rect -161 -142 -127 -108
rect 127 -142 161 -108
<< metal1 >>
rect -274 155 -208 160
rect -274 103 -268 155
rect -215 103 -208 155
rect -274 98 -208 103
rect -113 70 -79 280
rect 79 70 113 280
rect 207 155 273 160
rect 207 103 213 155
rect 266 103 273 155
rect 207 98 273 103
rect -321 64 -255 70
rect -321 -63 -311 64
rect -259 -63 -255 64
rect -321 -70 -255 -63
rect -225 64 -159 70
rect -225 -63 -215 64
rect -163 -63 -159 64
rect -225 -70 -159 -63
rect -119 58 -73 70
rect -119 -58 -113 58
rect -79 -58 -73 58
rect -119 -70 -73 -58
rect -33 64 33 70
rect -33 -63 -23 64
rect 29 -63 33 64
rect -33 -70 33 -63
rect 73 58 119 70
rect 73 -58 79 58
rect 113 -58 119 58
rect 73 -70 119 -58
rect 159 64 225 70
rect 159 -63 169 64
rect 221 -63 225 64
rect 159 -70 225 -63
rect 255 64 321 70
rect 255 -63 265 64
rect 317 -63 321 64
rect 255 -70 321 -63
rect -173 -108 -115 -102
rect 115 -108 173 -102
rect -305 -142 -161 -108
rect -127 -142 -111 -108
rect 115 -142 127 -108
rect 161 -142 305 -108
rect -173 -148 -115 -142
rect 115 -148 173 -142
<< via1 >>
rect -268 146 -215 155
rect -268 112 -258 146
rect -258 112 -224 146
rect -224 112 -215 146
rect -268 103 -215 112
rect 213 146 266 155
rect 213 112 223 146
rect 223 112 257 146
rect 257 112 266 146
rect 213 103 266 112
rect -311 58 -259 64
rect -311 -58 -305 58
rect -305 -58 -271 58
rect -271 -58 -259 58
rect -311 -63 -259 -58
rect -215 58 -163 64
rect -215 -58 -209 58
rect -209 -58 -175 58
rect -175 -58 -163 58
rect -215 -63 -163 -58
rect -23 58 29 64
rect -23 -58 -17 58
rect -17 -58 17 58
rect 17 -58 29 58
rect -23 -63 29 -58
rect 169 58 221 64
rect 169 -58 175 58
rect 175 -58 209 58
rect 209 -58 221 58
rect 169 -63 221 -58
rect 265 58 317 64
rect 265 -58 271 58
rect 271 -58 305 58
rect 305 -58 317 58
rect 265 -63 317 -58
<< metal2 >>
rect -37 173 37 182
rect -274 155 -208 160
rect -274 103 -268 155
rect -215 146 -208 155
rect -37 146 -28 173
rect -215 117 -28 146
rect 28 146 37 173
rect 207 155 273 160
rect 207 146 213 155
rect 28 117 213 146
rect -215 112 213 117
rect -215 103 -208 112
rect -274 98 -208 103
rect 207 103 213 112
rect 266 103 273 155
rect 207 98 273 103
rect -321 64 -255 70
rect -321 -63 -311 64
rect -259 17 -255 64
rect -225 64 -159 70
rect -225 17 -215 64
rect -259 -17 -215 17
rect -259 -63 -255 -17
rect -321 -70 -255 -63
rect -225 -63 -215 -17
rect -163 17 -159 64
rect -33 64 33 70
rect -33 17 -23 64
rect -163 -17 -23 17
rect -163 -63 -159 -17
rect -225 -70 -159 -63
rect -33 -63 -23 -17
rect 29 17 33 64
rect 159 64 225 70
rect 159 17 169 64
rect 29 -17 169 17
rect 29 -63 33 -17
rect -33 -70 33 -63
rect 159 -63 169 -17
rect 221 17 225 64
rect 255 64 321 70
rect 255 17 265 64
rect 221 -17 265 17
rect 221 -63 225 -17
rect 159 -70 225 -63
rect 255 -63 265 -17
rect 317 -63 321 64
rect 255 -70 321 -63
rect -22 -280 22 -70
<< via2 >>
rect -28 117 28 173
<< metal3 >>
rect -30 178 30 280
rect -33 173 33 178
rect -33 117 -28 173
rect 28 117 33 173
rect -33 112 33 117
<< properties >>
string FIXED_BBOX -402 -227 402 227
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.7 l 0.150 m 1 nf 6 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
