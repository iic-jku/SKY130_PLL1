magic
tech sky130A
magscale 1 2
timestamp 1663428559
<< metal1 >>
rect -237 353 -121 387
rect -63 353 4845 387
rect 5383 353 5755 387
rect 6677 353 6793 387
rect -237 -916 -203 353
rect 3138 302 3208 311
rect 3138 250 3147 302
rect 3199 250 3208 302
rect 3138 241 3208 250
rect 1371 119 1377 128
rect 1089 85 1377 119
rect 1371 76 1377 85
rect 1429 76 1435 128
rect 1481 76 1487 128
rect 1539 119 1545 128
rect 1539 85 1907 119
rect 1539 76 1545 85
rect -166 -182 -114 -176
rect -114 -225 -25 -191
rect 1089 -225 1907 -191
rect -166 -240 -114 -234
rect -63 -493 1127 -459
rect 1371 -769 1377 -760
rect 1089 -803 1377 -769
rect 1371 -812 1377 -803
rect 1429 -812 1435 -760
rect 1591 -769 1625 -225
rect 3156 -441 3190 241
rect 3232 76 3238 128
rect 3290 119 3296 128
rect 3290 85 3647 119
rect 3290 76 3296 85
rect 4595 -79 4601 -27
rect 4653 -79 4659 -27
rect 5537 -79 5543 -27
rect 5595 -79 5601 -27
rect 6759 -338 6793 353
rect 6741 -347 6811 -338
rect 6741 -399 6750 -347
rect 6802 -399 6811 -347
rect 6741 -408 6811 -399
rect 1869 -493 2867 -459
rect 3156 -475 4941 -441
rect 5287 -475 5947 -441
rect 3156 -659 3190 -475
rect 3147 -665 3199 -659
rect 3147 -723 3199 -717
rect 1591 -803 1907 -769
rect 2253 -803 3647 -769
rect 3147 -855 3199 -849
rect 3147 -913 3199 -907
rect -255 -925 -185 -916
rect -255 -977 -246 -925
rect -194 -977 -185 -925
rect -255 -986 -185 -977
rect 3156 -1019 3190 -913
rect 513 -1053 1127 -1019
rect 1185 -1053 3551 -1019
rect 3609 -1053 4031 -1019
rect 2303 -1329 2337 -1053
rect 3563 -1329 3597 -1053
rect 1869 -1363 2291 -1329
rect 3609 -1363 4031 -1329
rect 1481 -1622 1487 -1570
rect 1539 -1579 1545 -1570
rect 1539 -1613 1907 -1579
rect 1539 -1622 1545 -1613
rect 3232 -1622 3238 -1570
rect 3290 -1579 3296 -1570
rect 3290 -1613 3647 -1579
rect 3290 -1622 3296 -1613
<< via1 >>
rect 3147 250 3199 302
rect 1377 76 1429 128
rect 1487 76 1539 128
rect -166 -234 -114 -182
rect 1377 -812 1429 -760
rect 3238 76 3290 128
rect 4601 -79 4653 -27
rect 5543 -79 5595 -27
rect 6750 -399 6802 -347
rect 3147 -717 3199 -665
rect 3147 -907 3199 -855
rect -246 -977 -194 -925
rect 1487 -1622 1539 -1570
rect 3238 -1622 3290 -1570
<< metal2 >>
rect 3143 311 3203 315
rect 3138 306 3208 311
rect 3138 246 3143 306
rect 3203 246 3208 306
rect 3138 241 3208 246
rect 4797 304 4853 313
rect 6670 306 6726 315
rect 4853 254 4858 298
rect 3143 237 3203 241
rect 4797 239 4853 248
rect 5431 246 5708 306
rect 6665 256 6670 300
rect 6670 241 6726 250
rect -172 -191 -166 -182
rect -307 -225 -166 -191
rect -172 -234 -166 -225
rect -114 -234 -108 -182
rect 502 -272 562 166
rect 1377 128 1429 134
rect 1377 70 1429 76
rect 1487 128 1539 134
rect 1487 70 1539 76
rect 1386 -38 1420 70
rect 1376 -47 1432 -38
rect 1376 -112 1432 -103
rect 502 -492 562 -483
rect 502 -561 562 -552
rect 510 -609 554 -561
rect 510 -653 842 -609
rect 798 -842 842 -653
rect 1386 -754 1420 -112
rect 1496 -345 1530 70
rect 2338 -272 2398 166
rect 3238 128 3290 134
rect 3238 70 3290 76
rect 3247 -345 3281 70
rect 3792 -47 3848 -38
rect 3990 -53 4034 166
rect 4601 -27 4653 -21
rect 4595 -53 4601 -32
rect 3848 -79 4601 -53
rect 5543 -27 5595 -21
rect 5537 -74 5543 -32
rect 3848 -97 4653 -79
rect 5543 -85 5595 -79
rect 3792 -112 3848 -103
rect 1485 -354 1541 -345
rect 1485 -419 1541 -410
rect 3236 -354 3292 -345
rect 3236 -419 3292 -410
rect 1377 -760 1429 -754
rect 1377 -818 1429 -812
rect -250 -916 -190 -912
rect -255 -921 -185 -916
rect -255 -981 -250 -921
rect -190 -981 -185 -921
rect -255 -986 -185 -981
rect -250 -990 -190 -986
rect 1496 -1564 1530 -419
rect 3141 -717 3147 -665
rect 3199 -717 3205 -665
rect 3156 -855 3190 -717
rect 3141 -907 3147 -855
rect 3199 -907 3205 -855
rect 2058 -1401 2102 -981
rect 3247 -1564 3281 -419
rect 3798 -557 3842 -112
rect 4893 -345 4949 -336
rect 4949 -395 4954 -351
rect 4893 -410 4949 -401
rect 5335 -403 5899 -343
rect 6478 -345 6534 -336
rect 6746 -338 6806 -334
rect 6473 -395 6478 -351
rect 6478 -410 6534 -401
rect 6741 -343 6811 -338
rect 6741 -403 6746 -343
rect 6806 -403 6811 -343
rect 6741 -408 6811 -403
rect 6746 -412 6806 -408
rect 3790 -566 3850 -557
rect 3790 -635 3850 -626
rect 3798 -1401 3842 -981
rect 1487 -1570 1539 -1564
rect 1487 -1628 1539 -1622
rect 3238 -1570 3290 -1564
rect 3238 -1628 3290 -1622
<< via2 >>
rect 3143 302 3203 306
rect 3143 250 3147 302
rect 3147 250 3199 302
rect 3199 250 3203 302
rect 3143 246 3203 250
rect 4797 248 4853 304
rect 6670 250 6726 306
rect 1376 -103 1432 -47
rect 502 -552 562 -492
rect 3792 -103 3848 -47
rect 1485 -410 1541 -354
rect 3236 -410 3292 -354
rect -250 -925 -190 -921
rect -250 -977 -246 -925
rect -246 -977 -194 -925
rect -194 -977 -190 -925
rect -250 -981 -190 -977
rect 4893 -401 4949 -345
rect 6478 -401 6534 -345
rect 6746 -347 6806 -343
rect 6746 -399 6750 -347
rect 6750 -399 6802 -347
rect 6802 -399 6806 -347
rect 6746 -403 6806 -399
rect 3790 -626 3850 -566
<< metal3 >>
rect 3143 311 3203 315
rect 3138 306 3208 311
rect 4792 306 4858 309
rect -307 246 -177 306
rect 1241 246 1755 306
rect 2981 246 3143 306
rect 3203 246 3495 306
rect 4529 304 4858 306
rect 4529 248 4797 304
rect 4853 248 4858 304
rect 4529 246 4858 248
rect 3138 241 3208 246
rect 4792 243 4858 246
rect 6665 308 6731 311
rect 6665 306 6863 308
rect 6665 250 6670 306
rect 6726 250 6863 306
rect 6665 248 6863 250
rect 6665 245 6731 248
rect 3143 237 3203 241
rect 1371 -45 1437 -42
rect 3787 -45 3853 -42
rect 1371 -47 3853 -45
rect 1371 -103 1376 -47
rect 1432 -103 3792 -47
rect 3848 -103 3853 -47
rect 1371 -105 3853 -103
rect 1371 -108 1437 -105
rect 3787 -108 3853 -105
rect 6746 -338 6806 -334
rect 4888 -343 4954 -340
rect 4275 -345 4954 -343
rect 1480 -352 1546 -349
rect 3231 -352 3297 -349
rect 1241 -354 1546 -352
rect 1241 -410 1485 -354
rect 1541 -410 1546 -354
rect 1241 -412 1546 -410
rect 2981 -354 3297 -352
rect 2981 -410 3236 -354
rect 3292 -410 3297 -354
rect 2981 -412 3297 -410
rect 502 -487 562 -414
rect 1480 -415 1546 -412
rect 2309 -414 2427 -412
rect 497 -492 567 -487
rect 497 -552 502 -492
rect 562 -552 567 -492
rect 497 -557 567 -552
rect 2338 -601 2398 -414
rect 3231 -415 3297 -412
rect 4275 -401 4893 -345
rect 4949 -401 4954 -345
rect 4275 -403 4954 -401
rect 2050 -661 2398 -601
rect 3785 -566 3855 -561
rect 3785 -626 3790 -566
rect 3850 -626 3855 -566
rect 3785 -631 3855 -626
rect 2050 -839 2110 -661
rect 3790 -839 3850 -631
rect -250 -916 -190 -912
rect -255 -921 -185 -916
rect -307 -981 -250 -921
rect -190 -981 399 -921
rect 1241 -981 1431 -921
rect -255 -986 -185 -981
rect -250 -990 -190 -986
rect 1370 -1481 1430 -981
rect 4275 -1481 4335 -403
rect 4888 -406 4954 -403
rect 6473 -343 6539 -340
rect 6741 -343 6811 -338
rect 6473 -345 6746 -343
rect 6473 -401 6478 -345
rect 6534 -401 6746 -345
rect 6473 -403 6746 -401
rect 6806 -403 6863 -343
rect 6473 -406 6539 -403
rect 6741 -408 6811 -403
rect 6746 -412 6806 -408
rect 1370 -1541 1755 -1481
rect 2405 -1541 3495 -1481
rect 4145 -1541 4335 -1481
use simple2_inv  simple2_inv_0
timestamp 1661797765
transform 1 0 5611 0 1 0
box -42 -613 1252 525
use simple_inv  simple_inv_0
timestamp 1660926584
transform 1 0 4712 0 1 0
box -53 -613 857 525
use d_ff_n2  sky130_fd_pr__nfet_01v8_GVQ53W_0
timestamp 1663426905
transform 1 0 2080 0 1 -911
box -455 -280 455 280
use d_ff_n2  sky130_fd_pr__nfet_01v8_GVQ53W_1
timestamp 1663426905
transform -1 0 2080 0 -1 -1471
box -455 -280 455 280
use d_ff_n2  sky130_fd_pr__nfet_01v8_GVQ53W_2
timestamp 1663426905
transform 1 0 3820 0 1 -911
box -455 -280 455 280
use d_ff_n2  sky130_fd_pr__nfet_01v8_GVQ53W_3
timestamp 1663426905
transform -1 0 3820 0 -1 -1471
box -455 -280 455 280
use d_ff_n1  sky130_fd_pr__nfet_01v8_WWA63A_0
timestamp 1663426905
transform 1 0 820 0 1 -911
box -551 -280 551 280
use d_ff_p2  sky130_fd_pr__pfet_01v8_BD2UMN_0
timestamp 1663426905
transform 1 0 2368 0 1 236
box -743 -289 743 289
use d_ff_p2  sky130_fd_pr__pfet_01v8_BD2UMN_1
timestamp 1663426905
transform -1 0 2368 0 -1 -342
box -743 -289 743 289
use d_ff_p3  sky130_fd_pr__pfet_01v8_BDAGKN_0
timestamp 1663426905
transform 1 0 4012 0 1 236
box -647 -289 647 289
use d_ff_p1  sky130_fd_pr__pfet_01v8_BDS2ZN_0
timestamp 1663426905
transform 1 0 532 0 1 236
box -839 -289 839 289
use d_ff_p1  sky130_fd_pr__pfet_01v8_BDS2ZN_1
timestamp 1663426905
transform -1 0 532 0 -1 -342
box -839 -289 839 289
<< end >>
