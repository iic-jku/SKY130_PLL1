magic
tech sky130A
magscale 1 2
timestamp 1668153059
<< pwell >>
rect -2496 -2369 2460 2369
<< psubdiff >>
rect -2460 2299 -2364 2333
rect 2364 2299 2460 2333
rect -2460 2237 -2426 2299
rect 2426 2237 2460 2299
rect -2460 -2299 -2426 -2237
rect 2426 -2299 2460 -2237
rect -2460 -2333 -2364 -2299
rect 2364 -2333 2460 -2299
<< psubdiffcont >>
rect -2364 2299 2364 2333
rect -2460 -2237 -2426 2237
rect 2426 -2237 2460 2237
rect -2364 -2333 2364 -2299
<< xpolycontact >>
rect -2330 1771 -1760 2203
rect -2330 -2203 -1760 -1771
rect -1512 1771 -942 2203
rect -1512 -2203 -942 -1771
rect -694 1771 -124 2203
rect -694 -2203 -124 -1771
rect 124 1771 694 2203
rect 124 -2203 694 -1771
rect 942 1771 1512 2203
rect 942 -2203 1512 -1771
rect 1760 1771 2330 2203
rect 1760 -2203 2330 -1771
<< ppolyres >>
rect -2330 -1771 -1760 1771
rect -1512 -1771 -942 1771
rect -694 -1771 -124 1771
rect 124 -1771 694 1771
rect 942 -1771 1512 1771
rect 1760 -1771 2330 1771
<< locali >>
rect -2460 2299 -2364 2333
rect 2364 2299 2460 2333
rect -2460 2237 -2426 2299
rect 2426 2237 2460 2299
rect -2460 -2299 -2426 -2237
rect 2426 -2299 2460 -2237
rect -2460 -2333 -2364 -2299
rect 2364 -2333 2460 -2299
<< viali >>
rect -2314 1788 -1776 2185
rect -1496 1788 -958 2185
rect -678 1788 -140 2185
rect 140 1788 678 2185
rect 958 1788 1496 2185
rect 1776 1788 2314 2185
rect -2314 -2185 -1776 -1788
rect -1496 -2185 -958 -1788
rect -678 -2185 -140 -1788
rect 140 -2185 678 -1788
rect 958 -2185 1496 -1788
rect 1776 -2185 2314 -1788
<< metal1 >>
rect -2326 2185 -1764 2191
rect -2326 1788 -2314 2185
rect -1776 1788 -1764 2185
rect -2326 1782 -1764 1788
rect -1508 2185 -946 2191
rect -1508 1788 -1496 2185
rect -958 1788 -946 2185
rect -1508 1782 -946 1788
rect -694 2185 694 2206
rect -694 1788 -678 2185
rect -140 1788 140 2185
rect 678 1788 694 2185
rect -694 1772 694 1788
rect 946 2185 1508 2191
rect 946 1788 958 2185
rect 1496 1788 1508 2185
rect 946 1782 1508 1788
rect 1764 2185 2326 2191
rect 1764 1788 1776 2185
rect 2314 1788 2326 2185
rect 1764 1782 2326 1788
rect -2330 -1788 -1760 -1771
rect -2330 -2185 -2314 -1788
rect -1776 -2185 -1760 -1788
rect -2330 -2203 -1760 -2185
rect -1512 -1788 -124 -1770
rect -1512 -2185 -1496 -1788
rect -958 -2185 -678 -1788
rect -140 -2185 -124 -1788
rect -1512 -2204 -124 -2185
rect 124 -1788 1512 -1768
rect 124 -2185 140 -1788
rect 678 -2185 958 -1788
rect 1496 -2185 1512 -1788
rect 124 -2202 1512 -2185
rect 1760 -1788 2330 -1771
rect 1760 -2185 1776 -1788
rect 2314 -2185 2330 -1788
rect 1760 -2203 2330 -2185
<< via1 >>
rect -1496 1788 -958 2185
rect 958 1788 1496 2185
rect -2314 -2185 -1776 -1788
rect 1776 -2185 2314 -1788
<< metal2 >>
rect -1512 2185 -942 2830
rect -1512 1788 -1496 2185
rect -958 1788 -942 2185
rect -1512 1771 -942 1788
rect 942 2185 1512 2830
rect 942 1788 958 2185
rect 1496 1788 1512 2185
rect 942 1771 1512 1788
rect -2330 -1788 2330 -1771
rect -2330 -2185 -2314 -1788
rect -1776 -2185 1776 -1788
rect 2314 -2185 2330 -1788
rect -2330 -2203 2330 -2185
<< res2p85 >>
rect -2332 -1773 -1758 1773
rect -1514 -1773 -940 1773
rect -696 -1773 -122 1773
rect 122 -1773 696 1773
rect 940 -1773 1514 1773
rect 1758 -1773 2332 1773
<< properties >>
string FIXED_BBOX -2443 -2316 2443 2316
string gencell sky130_fd_pr__res_high_po_2p85
string library sky130
string parameters w 2.850 l 17.71 m 1 nx 6 wmin 2.850 lmin 0.50 rho 319.8 val 2.0k dummy 0 dw 0.0 term 19.188 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} full_metal 1 wmax 2.850 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
