magic
tech sky130A
timestamp 1654415419
<< pwell >>
rect -227 -140 227 140
<< nmos >>
rect -127 -35 -112 35
rect -79 -35 -64 35
rect -31 -35 -16 35
rect 16 -35 31 35
rect 64 -35 79 35
rect 112 -35 127 35
<< ndiff >>
rect -158 29 -127 35
rect -158 -29 -152 29
rect -135 -29 -127 29
rect -158 -35 -127 -29
rect -112 29 -79 35
rect -112 -29 -104 29
rect -87 -29 -79 29
rect -112 -35 -79 -29
rect -64 29 -31 35
rect -64 -29 -56 29
rect -39 -29 -31 29
rect -64 -35 -31 -29
rect -16 29 16 35
rect -16 -29 -8 29
rect 8 -29 16 29
rect -16 -35 16 -29
rect 31 29 64 35
rect 31 -29 39 29
rect 56 -29 64 29
rect 31 -35 64 -29
rect 79 29 112 35
rect 79 -29 87 29
rect 104 -29 112 29
rect 79 -35 112 -29
rect 127 29 158 35
rect 127 -29 135 29
rect 152 -29 158 29
rect 127 -35 158 -29
<< ndiffc >>
rect -152 -29 -135 29
rect -104 -29 -87 29
rect -56 -29 -39 29
rect -8 -29 8 29
rect 39 -29 56 29
rect 87 -29 104 29
rect 135 -29 152 29
<< psubdiff >>
rect -209 105 -161 122
rect 161 105 209 122
rect -209 74 -192 105
rect 192 74 209 105
rect -209 -105 -192 -74
rect 192 -105 209 -74
rect -209 -122 -161 -105
rect 161 -122 209 -105
<< psubdiffcont >>
rect -161 105 161 122
rect -209 -74 -192 74
rect 192 -74 209 74
rect -161 -122 161 -105
<< poly >>
rect -88 71 88 79
rect -88 54 -80 71
rect -63 54 -32 71
rect -15 54 15 71
rect 32 54 63 71
rect 80 54 88 71
rect -127 35 -112 48
rect -88 46 88 54
rect -79 35 -64 46
rect -31 35 -16 46
rect 16 35 31 46
rect 64 35 79 46
rect 112 35 127 48
rect -127 -51 -112 -35
rect -79 -48 -64 -35
rect -31 -48 -16 -35
rect 16 -48 31 -35
rect 64 -48 79 -35
rect 112 -51 127 -35
rect -136 -59 -103 -51
rect -136 -76 -128 -59
rect -111 -76 -103 -59
rect -136 -84 -103 -76
rect 103 -59 136 -51
rect 103 -76 111 -59
rect 128 -76 136 -59
rect 103 -84 136 -76
<< polycont >>
rect -80 54 -63 71
rect -32 54 -15 71
rect 15 54 32 71
rect 63 54 80 71
rect -128 -76 -111 -59
rect 111 -76 128 -59
<< locali >>
rect -209 105 -161 122
rect 161 105 209 122
rect -209 74 -192 105
rect 192 74 209 105
rect -88 54 -80 71
rect -63 54 -32 71
rect -15 54 15 71
rect 32 54 63 71
rect 80 54 88 71
rect -152 29 -135 37
rect -152 -37 -135 -29
rect -104 29 -87 37
rect -104 -37 -87 -29
rect -56 29 -39 37
rect -56 -37 -39 -29
rect -8 29 8 37
rect -8 -37 8 -29
rect 39 29 56 37
rect 39 -37 56 -29
rect 87 29 104 37
rect 87 -37 104 -29
rect 135 29 152 37
rect 135 -37 152 -29
rect -209 -105 -192 -74
rect -136 -76 -128 -59
rect -111 -76 -103 -59
rect 103 -76 111 -59
rect 128 -76 136 -59
rect 192 -105 209 -74
rect -209 -122 -161 -105
rect 161 -122 209 -105
<< viali >>
rect -80 54 -63 71
rect -32 54 -15 71
rect 15 54 32 71
rect 63 54 80 71
rect -152 -29 -135 29
rect -104 -29 -87 29
rect -56 -29 -39 29
rect -8 -29 8 29
rect 39 -29 56 29
rect 87 -29 104 29
rect 135 -29 152 29
rect -128 -76 -111 -59
rect 111 -76 128 -59
<< metal1 >>
rect -86 71 -57 74
rect -38 71 -9 74
rect 9 71 38 74
rect 57 71 86 74
rect -86 54 -80 71
rect -63 54 -32 71
rect -15 54 15 71
rect 32 54 63 71
rect 80 54 86 71
rect -86 51 -57 54
rect -38 51 -9 54
rect 9 51 38 54
rect 57 51 86 54
rect -155 29 -132 35
rect -155 -29 -152 29
rect -135 -29 -132 29
rect -155 -35 -132 -29
rect -112 29 -79 35
rect -112 -29 -109 29
rect -83 -29 -79 29
rect -112 -35 -79 -29
rect -59 29 -36 35
rect -59 -29 -56 29
rect -39 -29 -36 29
rect -59 -35 -36 -29
rect -16 29 16 35
rect -16 -29 -13 29
rect 13 -29 16 29
rect -16 -35 16 -29
rect 36 29 59 35
rect 36 -29 39 29
rect 56 -29 59 29
rect 36 -35 59 -29
rect 79 29 112 35
rect 79 -29 82 29
rect 109 -29 112 29
rect 79 -35 112 -29
rect 132 29 155 35
rect 132 -29 135 29
rect 152 -29 155 29
rect 132 -35 155 -29
rect -136 -55 -103 -51
rect -136 -81 -133 -55
rect -107 -81 -103 -55
rect -136 -84 -103 -81
rect 103 -55 136 -51
rect 103 -81 107 -55
rect 133 -81 136 -55
rect 103 -84 136 -81
<< via1 >>
rect -109 -29 -104 29
rect -104 -29 -87 29
rect -87 -29 -83 29
rect -13 -29 -8 29
rect -8 -29 8 29
rect 8 -29 13 29
rect 82 -29 87 29
rect 87 -29 104 29
rect 104 -29 109 29
rect -133 -59 -107 -55
rect -133 -76 -128 -59
rect -128 -76 -111 -59
rect -111 -76 -107 -59
rect -133 -81 -107 -76
rect 107 -59 133 -55
rect 107 -76 111 -59
rect 111 -76 128 -59
rect 128 -76 133 -59
rect 107 -81 133 -76
<< metal2 >>
rect -112 29 -79 35
rect -112 -29 -109 29
rect -83 -18 -79 29
rect -16 29 16 35
rect -16 -18 -13 29
rect -83 -29 -13 -18
rect 13 -18 16 29
rect 79 29 112 35
rect 79 -18 82 29
rect 13 -29 82 -18
rect 109 -29 112 29
rect -112 -35 112 -29
rect -139 -53 -101 -49
rect -139 -82 -134 -53
rect -105 -82 -101 -53
rect -139 -87 -101 -82
rect -8 -140 8 -35
rect 101 -53 139 -49
rect 101 -82 105 -53
rect 134 -82 139 -53
rect 101 -87 139 -82
<< via2 >>
rect -134 -55 -105 -53
rect -134 -81 -133 -55
rect -133 -81 -107 -55
rect -107 -81 -105 -55
rect -134 -82 -105 -81
rect 105 -55 134 -53
rect 105 -81 107 -55
rect 107 -81 133 -55
rect 133 -81 134 -55
rect 105 -82 134 -81
<< metal3 >>
rect -139 -53 -101 -49
rect 101 -53 139 -49
rect -139 -53 139 -53
rect -139 -82 -134 -53
rect -105 -82 105 -53
rect 134 -82 139 -53
rect -139 -83 139 -82
rect -139 -87 -101 -83
rect 101 -87 139 -83
<< properties >>
string FIXED_BBOX -201 -113 201 113
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.7 l 0.150 m 1 nf 6 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
