magic
tech sky130A
magscale 1 2
timestamp 1654967793
<< nwell >>
rect -743 -289 743 289
<< pmos >>
rect -543 -70 -513 70
rect -447 -70 -417 70
rect -351 -70 -321 70
rect -255 -70 -225 70
rect -159 -70 -129 70
rect -63 -70 -33 70
rect 33 -70 63 70
rect 129 -70 159 70
rect 225 -70 255 70
rect 321 -70 351 70
rect 417 -70 447 70
rect 513 -70 543 70
<< pdiff >>
rect -605 58 -543 70
rect -605 -58 -593 58
rect -559 -58 -543 58
rect -605 -70 -543 -58
rect -513 58 -447 70
rect -513 -58 -497 58
rect -463 -58 -447 58
rect -513 -70 -447 -58
rect -417 58 -351 70
rect -417 -58 -401 58
rect -367 -58 -351 58
rect -417 -70 -351 -58
rect -321 58 -255 70
rect -321 -58 -305 58
rect -271 -58 -255 58
rect -321 -70 -255 -58
rect -225 58 -159 70
rect -225 -58 -209 58
rect -175 -58 -159 58
rect -225 -70 -159 -58
rect -129 58 -63 70
rect -129 -58 -113 58
rect -79 -58 -63 58
rect -129 -70 -63 -58
rect -33 58 33 70
rect -33 -58 -17 58
rect 17 -58 33 58
rect -33 -70 33 -58
rect 63 58 129 70
rect 63 -58 79 58
rect 113 -58 129 58
rect 63 -70 129 -58
rect 159 58 225 70
rect 159 -58 175 58
rect 209 -58 225 58
rect 159 -70 225 -58
rect 255 58 321 70
rect 255 -58 271 58
rect 305 -58 321 58
rect 255 -70 321 -58
rect 351 58 417 70
rect 351 -58 367 58
rect 401 -58 417 58
rect 351 -70 417 -58
rect 447 58 513 70
rect 447 -58 463 58
rect 497 -58 513 58
rect 447 -70 513 -58
rect 543 58 605 70
rect 543 -58 559 58
rect 593 -58 605 58
rect 543 -70 605 -58
<< pdiffc >>
rect -593 -58 -559 58
rect -497 -58 -463 58
rect -401 -58 -367 58
rect -305 -58 -271 58
rect -209 -58 -175 58
rect -113 -58 -79 58
rect -17 -58 17 58
rect 79 -58 113 58
rect 175 -58 209 58
rect 271 -58 305 58
rect 367 -58 401 58
rect 463 -58 497 58
rect 559 -58 593 58
<< nsubdiff >>
rect -707 219 -611 253
rect 611 219 707 253
rect -707 157 -673 219
rect 673 157 707 219
rect -707 -219 -673 -157
rect 673 -219 707 -157
rect -707 -253 -611 -219
rect 611 -253 707 -219
<< nsubdiffcont >>
rect -611 219 611 253
rect -707 -157 -673 157
rect 673 -157 707 157
rect -611 -253 611 -219
<< poly >>
rect -465 151 465 167
rect -465 117 -449 151
rect -415 117 -353 151
rect -319 117 -257 151
rect -223 117 -161 151
rect -127 117 -65 151
rect -31 117 31 151
rect 65 117 127 151
rect 161 117 223 151
rect 257 117 319 151
rect 353 117 415 151
rect 449 117 465 151
rect -465 101 465 117
rect -543 70 -513 96
rect -447 70 -417 101
rect -351 70 -321 101
rect -255 70 -225 101
rect -159 70 -129 101
rect -63 70 -33 101
rect 33 70 63 101
rect 129 70 159 101
rect 225 70 255 101
rect 321 70 351 101
rect 417 70 447 101
rect 513 70 543 96
rect -543 -101 -513 -70
rect -447 -96 -417 -70
rect -351 -96 -321 -70
rect -255 -96 -225 -70
rect -159 -96 -129 -70
rect -63 -96 -33 -70
rect 33 -96 63 -70
rect 129 -96 159 -70
rect 225 -96 255 -70
rect 321 -96 351 -70
rect 417 -96 447 -70
rect 513 -101 543 -70
rect -561 -117 -495 -101
rect -561 -151 -545 -117
rect -511 -151 -495 -117
rect -561 -167 -495 -151
rect 495 -117 561 -101
rect 495 -151 511 -117
rect 545 -151 561 -117
rect 495 -167 561 -151
<< polycont >>
rect -449 117 -415 151
rect -353 117 -319 151
rect -257 117 -223 151
rect -161 117 -127 151
rect -65 117 -31 151
rect 31 117 65 151
rect 127 117 161 151
rect 223 117 257 151
rect 319 117 353 151
rect 415 117 449 151
rect -545 -151 -511 -117
rect 511 -151 545 -117
<< locali >>
rect -707 219 -611 253
rect 611 219 707 253
rect -707 157 -673 219
rect 673 157 707 219
rect -465 117 -449 151
rect -415 117 -353 151
rect -319 117 -257 151
rect -223 117 -161 151
rect -127 117 -65 151
rect -31 117 31 151
rect 65 117 127 151
rect 161 117 223 151
rect 257 117 319 151
rect 353 117 415 151
rect 449 117 465 151
rect -593 58 -559 74
rect -593 -74 -559 -58
rect -497 58 -463 74
rect -497 -74 -463 -58
rect -401 58 -367 74
rect -401 -74 -367 -58
rect -305 58 -271 74
rect -305 -74 -271 -58
rect -209 58 -175 74
rect -209 -74 -175 -58
rect -113 58 -79 74
rect -113 -74 -79 -58
rect -17 58 17 74
rect -17 -74 17 -58
rect 79 58 113 74
rect 79 -74 113 -58
rect 175 58 209 74
rect 175 -74 209 -58
rect 271 58 305 74
rect 271 -74 305 -58
rect 367 58 401 74
rect 367 -74 401 -58
rect 463 58 497 74
rect 463 -74 497 -58
rect 559 58 593 74
rect 559 -74 593 -58
rect -561 -151 -545 -117
rect -511 -151 -495 -117
rect 495 -151 511 -117
rect 545 -151 561 -117
rect -707 -219 -673 -157
rect 673 -219 707 -157
rect -707 -253 -611 -219
rect 611 -253 707 -219
<< viali >>
rect -449 117 -415 151
rect -353 117 -319 151
rect -257 117 -223 151
rect -161 117 -127 151
rect -65 117 -31 151
rect 31 117 65 151
rect 127 117 161 151
rect 223 117 257 151
rect 319 117 353 151
rect 415 117 449 151
rect -593 -58 -559 58
rect -497 -58 -463 58
rect -401 -58 -367 58
rect -305 -58 -271 58
rect -209 -58 -175 58
rect -113 -58 -79 58
rect -17 -58 17 58
rect 79 -58 113 58
rect 175 -58 209 58
rect 271 -58 305 58
rect 367 -58 401 58
rect 463 -58 497 58
rect 559 -58 593 58
rect -545 -151 -511 -117
rect 511 -151 545 -117
<< metal1 >>
rect -272 160 -208 166
rect -461 151 -403 157
rect -365 151 -307 157
rect -272 151 -266 160
rect -214 151 -208 160
rect -173 151 -115 157
rect -77 151 -19 157
rect 19 151 77 157
rect 115 151 173 157
rect 211 151 269 157
rect 307 151 365 157
rect 403 151 461 157
rect -465 117 -449 151
rect -415 117 -353 151
rect -319 117 -266 151
rect -214 117 -161 151
rect -127 117 -65 151
rect -31 117 31 151
rect 65 117 127 151
rect 161 117 223 151
rect 257 117 319 151
rect 353 117 415 151
rect 449 117 465 151
rect -461 111 -403 117
rect -365 111 -307 117
rect -272 108 -266 117
rect -214 108 -208 117
rect -173 111 -115 117
rect -77 111 -19 117
rect 19 111 77 117
rect 115 111 173 117
rect 211 111 269 117
rect 307 111 365 117
rect 403 111 461 117
rect -272 102 -208 108
rect -599 58 -553 70
rect -599 -6 -593 58
rect -608 -14 -593 -6
rect -559 -6 -553 58
rect -512 64 -448 70
rect -512 12 -506 64
rect -454 12 -448 64
rect -512 6 -497 12
rect -559 -14 -544 -6
rect -608 -66 -602 -14
rect -550 -66 -544 -14
rect -608 -70 -544 -66
rect -503 -58 -497 6
rect -463 6 -448 12
rect -407 58 -361 70
rect -463 -58 -457 6
rect -407 -6 -401 58
rect -503 -70 -457 -58
rect -416 -14 -401 -6
rect -367 -6 -361 58
rect -320 64 -256 70
rect -320 12 -314 64
rect -262 12 -256 64
rect -320 6 -305 12
rect -367 -14 -352 -6
rect -416 -66 -410 -14
rect -358 -66 -352 -14
rect -416 -70 -352 -66
rect -311 -58 -305 6
rect -271 6 -256 12
rect -215 58 -169 70
rect -271 -58 -265 6
rect -215 -6 -209 58
rect -311 -70 -265 -58
rect -224 -14 -209 -6
rect -175 -6 -169 58
rect -128 64 -64 70
rect -128 12 -122 64
rect -70 12 -64 64
rect -128 6 -113 12
rect -175 -14 -160 -6
rect -224 -66 -218 -14
rect -166 -66 -160 -14
rect -224 -70 -160 -66
rect -119 -58 -113 6
rect -79 6 -64 12
rect -23 58 23 70
rect -79 -58 -73 6
rect -23 -6 -17 58
rect -119 -70 -73 -58
rect -32 -14 -17 -6
rect 17 -6 23 58
rect 64 64 128 70
rect 64 12 70 64
rect 122 12 128 64
rect 64 6 79 12
rect 17 -14 32 -6
rect -32 -66 -26 -14
rect 26 -66 32 -14
rect -32 -70 32 -66
rect 73 -58 79 6
rect 113 6 128 12
rect 169 58 215 70
rect 113 -58 119 6
rect 169 -6 175 58
rect 73 -70 119 -58
rect 160 -14 175 -6
rect 209 -6 215 58
rect 256 64 320 70
rect 256 12 262 64
rect 314 12 320 64
rect 256 6 271 12
rect 209 -14 224 -6
rect 160 -66 166 -14
rect 218 -66 224 -14
rect 160 -70 224 -66
rect 265 -58 271 6
rect 305 6 320 12
rect 361 58 407 70
rect 305 -58 311 6
rect 361 -6 367 58
rect 265 -70 311 -58
rect 352 -14 367 -6
rect 401 -6 407 58
rect 448 64 512 70
rect 448 12 454 64
rect 506 12 512 64
rect 448 6 463 12
rect 401 -14 416 -6
rect 352 -66 358 -14
rect 410 -66 416 -14
rect 352 -70 416 -66
rect 457 -58 463 6
rect 497 6 512 12
rect 553 58 599 70
rect 497 -58 503 6
rect 553 -6 559 58
rect 457 -70 503 -58
rect 544 -14 559 -6
rect 593 -6 599 58
rect 593 -14 608 -6
rect 544 -66 550 -14
rect 602 -66 608 -14
rect 544 -70 608 -66
rect -557 -117 -499 -111
rect 499 -117 557 -111
rect -557 -151 -545 -117
rect -511 -151 511 -117
rect 545 -151 557 -117
rect -557 -157 -499 -151
rect 499 -157 557 -151
<< via1 >>
rect -266 151 -214 160
rect -266 117 -257 151
rect -257 117 -223 151
rect -223 117 -214 151
rect -266 108 -214 117
rect -506 58 -454 64
rect -506 12 -497 58
rect -497 12 -463 58
rect -463 12 -454 58
rect -602 -58 -593 -14
rect -593 -58 -559 -14
rect -559 -58 -550 -14
rect -602 -66 -550 -58
rect -314 58 -262 64
rect -314 12 -305 58
rect -305 12 -271 58
rect -271 12 -262 58
rect -410 -58 -401 -14
rect -401 -58 -367 -14
rect -367 -58 -358 -14
rect -410 -66 -358 -58
rect -122 58 -70 64
rect -122 12 -113 58
rect -113 12 -79 58
rect -79 12 -70 58
rect -218 -58 -209 -14
rect -209 -58 -175 -14
rect -175 -58 -166 -14
rect -218 -66 -166 -58
rect 70 58 122 64
rect 70 12 79 58
rect 79 12 113 58
rect 113 12 122 58
rect -26 -58 -17 -14
rect -17 -58 17 -14
rect 17 -58 26 -14
rect -26 -66 26 -58
rect 262 58 314 64
rect 262 12 271 58
rect 271 12 305 58
rect 305 12 314 58
rect 166 -58 175 -14
rect 175 -58 209 -14
rect 209 -58 218 -14
rect 166 -66 218 -58
rect 454 58 506 64
rect 454 12 463 58
rect 463 12 497 58
rect 497 12 506 58
rect 358 -58 367 -14
rect 367 -58 401 -14
rect 401 -58 410 -14
rect 358 -66 410 -58
rect 550 -58 559 -14
rect 559 -58 593 -14
rect 593 -58 602 -14
rect 550 -66 602 -58
<< metal2 >>
rect -257 166 -223 289
rect -272 160 -208 166
rect -272 108 -266 160
rect -214 108 -208 160
rect -272 102 -208 108
rect -512 64 743 70
rect -512 12 -506 64
rect -454 36 -314 64
rect -454 12 -448 36
rect -512 6 -448 12
rect -320 12 -314 36
rect -262 36 -122 64
rect -262 12 -256 36
rect -320 6 -256 12
rect -128 12 -122 36
rect -70 36 70 64
rect -70 12 -64 36
rect -128 6 -64 12
rect 64 12 70 36
rect 122 36 262 64
rect 122 12 128 36
rect 64 6 128 12
rect 256 12 262 36
rect 314 36 454 64
rect 314 12 320 36
rect 256 6 320 12
rect 448 12 454 36
rect 506 36 743 64
rect 506 12 512 36
rect 448 6 512 12
rect -613 -12 -539 -3
rect -613 -68 -604 -12
rect -548 -68 -539 -12
rect -613 -77 -539 -68
rect -421 -12 -347 -3
rect -421 -68 -412 -12
rect -356 -68 -347 -12
rect -421 -77 -347 -68
rect -229 -12 -155 -3
rect -229 -68 -220 -12
rect -164 -68 -155 -12
rect -229 -77 -155 -68
rect -37 -12 37 -3
rect -37 -68 -28 -12
rect 28 -68 37 -12
rect -37 -77 37 -68
rect 155 -12 229 -3
rect 155 -68 164 -12
rect 220 -68 229 -12
rect 155 -77 229 -68
rect 347 -12 421 -3
rect 347 -68 356 -12
rect 412 -68 421 -12
rect 347 -77 421 -68
rect 539 -12 613 -3
rect 539 -68 548 -12
rect 604 -68 613 -12
rect 539 -77 613 -68
<< via2 >>
rect -604 -14 -548 -12
rect -604 -66 -602 -14
rect -602 -66 -550 -14
rect -550 -66 -548 -14
rect -604 -68 -548 -66
rect -412 -14 -356 -12
rect -412 -66 -410 -14
rect -410 -66 -358 -14
rect -358 -66 -356 -14
rect -412 -68 -356 -66
rect -220 -14 -164 -12
rect -220 -66 -218 -14
rect -218 -66 -166 -14
rect -166 -66 -164 -14
rect -220 -68 -164 -66
rect -28 -14 28 -12
rect -28 -66 -26 -14
rect -26 -66 26 -14
rect 26 -66 28 -14
rect -28 -68 28 -66
rect 164 -14 220 -12
rect 164 -66 166 -14
rect 166 -66 218 -14
rect 218 -66 220 -14
rect 164 -68 220 -66
rect 356 -14 412 -12
rect 356 -66 358 -14
rect 358 -66 410 -14
rect 410 -66 412 -14
rect 356 -68 412 -66
rect 548 -14 604 -12
rect 548 -66 550 -14
rect 550 -66 602 -14
rect 602 -66 604 -14
rect 548 -68 604 -66
<< metal3 >>
rect -613 -10 -539 -3
rect -421 -10 -347 -3
rect -229 -10 -155 -3
rect -37 -10 37 -3
rect 155 -10 229 -3
rect 347 -10 421 -3
rect 539 -10 613 -3
rect -613 -12 613 -10
rect -613 -68 -604 -12
rect -548 -68 -412 -12
rect -356 -68 -220 -12
rect -164 -68 -28 -12
rect 28 -68 164 -12
rect 220 -68 356 -12
rect 412 -68 548 -12
rect 604 -68 613 -12
rect -613 -70 613 -68
rect -613 -77 -539 -70
rect -421 -77 -347 -70
rect -229 -77 -155 -70
rect -37 -77 37 -70
rect 155 -77 229 -70
rect 347 -77 421 -70
rect 539 -77 613 -70
<< properties >>
string FIXED_BBOX -690 -236 690 236
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.7 l 0.15 m 1 nf 12 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
