magic
tech sky130A
magscale 1 2
timestamp 1668357910
<< nwell >>
rect 1079 4318 1270 4896
rect 4253 3700 4831 3817
<< metal1 >>
rect 4039 5308 4045 5313
rect 3806 5266 4045 5308
rect 4039 5261 4045 5266
rect 4097 5261 4103 5313
rect 5351 5260 5357 5312
rect 5409 5260 6386 5312
rect 4429 4619 4435 4677
rect 4493 4619 4812 4677
rect 4870 4619 4876 4677
rect 1222 4344 1274 4350
rect -1125 4297 -1029 4339
rect 1222 4286 1274 4292
rect 4128 3864 4180 3870
rect 4180 3817 4682 3859
rect 4128 3806 4180 3812
rect 6334 3318 6386 5260
rect 4200 3154 4206 3206
rect 4258 3154 4264 3206
rect 6334 3164 6511 3318
rect 6086 2524 6132 2579
rect 4107 2251 4113 2256
rect 3874 2209 4113 2251
rect 4107 2204 4113 2209
rect 4165 2204 4171 2256
rect 5569 2204 5575 2256
rect 5627 2251 5633 2256
rect 6208 2251 6214 2256
rect 5627 2209 6214 2251
rect 5627 2204 5633 2209
rect 6208 2204 6214 2209
rect 6266 2204 6272 2256
rect 6334 2160 6386 3164
rect 6468 2262 6510 2416
rect 6458 2256 6510 2262
rect 6458 2198 6510 2204
rect 6334 2108 6629 2160
<< via1 >>
rect 4045 5261 4097 5313
rect 5357 5260 5409 5312
rect 4435 4619 4493 4677
rect 4812 4619 4870 4677
rect 1222 4292 1274 4344
rect 4128 3812 4180 3864
rect 4206 3154 4258 3206
rect 4113 2204 4165 2256
rect 5575 2204 5627 2256
rect 6214 2204 6266 2256
rect 6458 2204 6510 2256
<< metal2 >>
rect 6153 5420 7253 5490
rect 4045 5313 4097 5319
rect 5357 5312 5409 5318
rect 4097 5266 4211 5308
rect 5239 5266 5357 5308
rect 4045 5255 4097 5261
rect 5357 5254 5409 5260
rect 4435 4677 4493 4683
rect 942 4607 1196 4677
rect 4005 4619 4435 4677
rect 4435 4613 4493 4619
rect 4812 4677 4870 4683
rect 6153 4677 6211 5420
rect 4870 4619 6211 4677
rect 4812 4613 4870 4619
rect 1126 4508 1196 4607
rect 4950 4589 5020 4619
rect 1126 4438 1698 4508
rect 1216 4339 1222 4344
rect 1037 4297 1222 4339
rect 1216 4292 1222 4297
rect 1274 4292 1280 4344
rect 3999 4297 4175 4339
rect 750 3968 1130 4038
rect 4133 3864 4175 4297
rect 4122 3812 4128 3864
rect 4180 3812 4186 3864
rect 4311 3793 4381 4050
rect 4311 3723 5704 3793
rect 3861 3469 4472 3539
rect 5111 3466 5181 3723
rect 4206 3206 4258 3212
rect 3999 3159 4206 3201
rect 4206 3148 4258 3154
rect 3993 1594 4063 2889
rect 4113 2256 4165 2262
rect 5575 2256 5627 2262
rect 4165 2209 4253 2251
rect 5304 2223 5575 2251
rect 5293 2209 5575 2223
rect 4113 2198 4165 2204
rect 5293 1873 5433 2209
rect 5575 2198 5627 2204
rect 6214 2256 6266 2262
rect 6452 2251 6458 2256
rect 6266 2209 6458 2251
rect 6452 2204 6458 2209
rect 6510 2204 6516 2256
rect 6214 2198 6266 2204
rect 5293 1724 5433 1733
rect 3984 1524 3993 1594
rect 4063 1524 4072 1594
rect 3993 1514 4063 1524
rect 5578 1356 5587 1594
rect 5657 1356 5774 1594
<< via2 >>
rect 5293 1733 5433 1873
rect 3993 1524 4063 1594
rect 5587 1356 5657 1594
<< metal3 >>
rect 5288 1873 5438 1878
rect 5288 1868 5293 1873
rect 5433 1868 5438 1873
rect 5288 1722 5438 1728
rect 3988 1594 4068 1599
rect 5582 1594 5662 1599
rect 3988 1524 3993 1594
rect 4063 1524 4342 1594
rect 3988 1519 4068 1524
rect 5474 1356 5587 1594
rect 5657 1356 5662 1594
rect 5474 1351 5662 1356
<< via3 >>
rect 5288 1733 5293 1868
rect 5293 1733 5433 1868
rect 5433 1733 5438 1868
rect 5288 1728 5438 1733
<< metal4 >>
rect 5293 1869 5433 1873
rect 5287 1868 5439 1869
rect 5287 1728 5288 1868
rect 5438 1728 5439 1868
rect 5287 1727 5439 1728
rect 5293 1494 5433 1727
use cap50f  cap50f_0
timestamp 1668357910
transform 1 0 4983 0 1 994
box -650 -600 550 600
use differential  differential_0
timestamp 1668357910
transform 1 0 1268 0 1 2620
box -145 0 2794 2276
use inv_buffer2  inv_buffer2_0
timestamp 1668357910
transform 1 0 -1125 0 1 3758
box 0 0 2204 1138
use ota_2  ota_2_0
timestamp 1668357910
transform 0 1 6334 -1 0 5490
box 0 -630 5276 1138
use tgate_1  tgate_1_0
timestamp 1668357910
transform 1 0 4472 0 -1 2790
box -261 -952 919 1138
use tgate_1  tgate_1_1
timestamp 1668357910
transform -1 0 5020 0 1 4727
box -261 -952 919 1138
<< labels >>
rlabel metal1 -1125 4297 -1029 4339 7 ref_in
port 1 n
rlabel metal1 3874 2209 3970 2251 0 vco_in
port 2 n
rlabel metal1 6086 2524 6132 2579 0 vbias
port 4 n
rlabel metal2 7183 5420 7253 5490 0 vdd
port 5 n
rlabel metal2 5704 1356 5774 1426 0 vss
port 6 n
rlabel metal2 4062 4619 4211 4677 5 vdd
rlabel metal1 3806 5266 3902 5308 7 v_out
port 3 n
<< end >>
