magic
tech sky130A
magscale 1 2
timestamp 1660729001
<< error_p >>
rect 307 151 365 157
rect 307 117 319 151
rect 307 111 365 117
rect -365 -117 -307 -111
rect -365 -151 -353 -117
rect -365 -157 -307 -151
<< nwell >>
rect -551 -289 551 289
<< pmos >>
rect -351 -70 -321 70
rect -255 -70 -225 70
rect -159 -70 -129 70
rect -63 -70 -33 70
rect 33 -70 63 70
rect 129 -70 159 70
rect 225 -70 255 70
rect 321 -70 351 70
<< pdiff >>
rect -417 58 -351 70
rect -417 -58 -401 58
rect -367 -58 -351 58
rect -417 -70 -351 -58
rect -321 58 -255 70
rect -321 -58 -305 58
rect -271 -58 -255 58
rect -321 -70 -255 -58
rect -225 58 -159 70
rect -225 -58 -209 58
rect -175 -58 -159 58
rect -225 -70 -159 -58
rect -129 58 -63 70
rect -129 -58 -113 58
rect -79 -58 -63 58
rect -129 -70 -63 -58
rect -33 58 33 70
rect -33 -58 -17 58
rect 17 -58 33 58
rect -33 -70 33 -58
rect 63 58 129 70
rect 63 -58 79 58
rect 113 -58 129 58
rect 63 -70 129 -58
rect 159 58 225 70
rect 159 -58 175 58
rect 209 -58 225 58
rect 159 -70 225 -58
rect 255 58 321 70
rect 255 -58 271 58
rect 305 -58 321 58
rect 255 -70 321 -58
rect 351 58 417 70
rect 351 -58 367 58
rect 401 -58 417 58
rect 351 -70 417 -58
<< pdiffc >>
rect -401 -58 -367 58
rect -305 -58 -271 58
rect -209 -58 -175 58
rect -113 -58 -79 58
rect -17 -58 17 58
rect 79 -58 113 58
rect 175 -58 209 58
rect 271 -58 305 58
rect 367 -58 401 58
<< nsubdiff >>
rect -515 219 -419 253
rect 419 219 515 253
rect -515 157 -481 219
rect 481 157 515 219
rect -515 -219 -481 -157
rect 481 -219 515 -157
rect -515 -253 -419 -219
rect 419 -253 515 -219
<< nsubdiffcont >>
rect -419 219 419 253
rect -515 -157 -481 157
rect 481 -157 515 157
rect -419 -253 419 -219
<< poly >>
rect -273 151 -207 167
rect -273 117 -257 151
rect -223 117 -207 151
rect -273 101 -207 117
rect -81 151 -15 167
rect -81 117 -65 151
rect -31 117 -15 151
rect -81 101 -15 117
rect 111 151 177 167
rect 111 117 127 151
rect 161 117 177 151
rect 111 101 177 117
rect 303 151 369 167
rect 303 117 319 151
rect 353 117 369 151
rect 303 101 369 117
rect -351 70 -321 96
rect -255 70 -225 101
rect -159 70 -129 96
rect -63 70 -33 101
rect 33 70 63 96
rect 129 70 159 101
rect 225 70 255 96
rect 321 70 351 101
rect -351 -101 -321 -70
rect -255 -96 -225 -70
rect -159 -101 -129 -70
rect -63 -96 -33 -70
rect 33 -101 63 -70
rect 129 -96 159 -70
rect 225 -101 255 -70
rect 321 -96 351 -70
rect -369 -117 -303 -101
rect -369 -151 -353 -117
rect -319 -151 -303 -117
rect -369 -167 -303 -151
rect -177 -117 -111 -101
rect -177 -151 -161 -117
rect -127 -151 -111 -117
rect -177 -167 -111 -151
rect 15 -117 81 -101
rect 15 -151 31 -117
rect 65 -151 81 -117
rect 15 -167 81 -151
rect 207 -117 273 -101
rect 207 -151 223 -117
rect 257 -151 273 -117
rect 207 -167 273 -151
<< polycont >>
rect -257 117 -223 151
rect -65 117 -31 151
rect 127 117 161 151
rect 319 117 353 151
rect -353 -151 -319 -117
rect -161 -151 -127 -117
rect 31 -151 65 -117
rect 223 -151 257 -117
<< locali >>
rect -515 219 -419 253
rect 419 219 515 253
rect -515 157 -481 219
rect 481 157 515 219
rect -273 117 -257 151
rect -223 117 -207 151
rect -81 117 -65 151
rect -31 117 -15 151
rect 111 117 127 151
rect 161 117 177 151
rect 303 117 319 151
rect 353 117 369 151
rect -401 58 -367 74
rect -401 -74 -367 -58
rect -305 58 -271 74
rect -305 -74 -271 -58
rect -209 58 -175 74
rect -209 -74 -175 -58
rect -113 58 -79 74
rect -113 -74 -79 -58
rect -17 58 17 74
rect -17 -74 17 -58
rect 79 58 113 74
rect 79 -74 113 -58
rect 175 58 209 74
rect 175 -74 209 -58
rect 271 58 305 74
rect 271 -74 305 -58
rect 367 58 401 74
rect 367 -74 401 -58
rect -369 -151 -353 -117
rect -319 -151 -303 -117
rect -177 -151 -161 -117
rect -127 -151 -111 -117
rect 15 -151 31 -117
rect 65 -151 81 -117
rect 207 -151 223 -117
rect 257 -151 273 -117
rect -515 -219 -481 -157
rect 481 -219 515 -157
rect -515 -253 -419 -219
rect 419 -253 515 -219
<< viali >>
rect -257 117 -223 151
rect -65 117 -31 151
rect 127 117 161 151
rect 319 117 353 151
rect -401 -58 -367 58
rect -305 -58 -271 58
rect -209 -58 -175 58
rect -113 -58 -79 58
rect -17 -58 17 58
rect 79 -58 113 58
rect 175 -58 209 58
rect 271 -58 305 58
rect 367 -58 401 58
rect -353 -151 -319 -117
rect -161 -151 -127 -117
rect 31 -151 65 -117
rect 223 -151 257 -117
<< metal1 >>
rect -362 160 -310 166
rect -269 151 -211 157
rect -310 117 -257 151
rect -223 117 -211 151
rect -269 111 -211 117
rect -77 151 -19 157
rect 115 151 173 157
rect -77 117 -65 151
rect -31 117 127 151
rect 161 117 173 151
rect -77 111 -19 117
rect 79 111 173 117
rect 307 151 365 157
rect 307 117 319 151
rect 353 117 365 151
rect 307 111 365 117
rect -362 102 -310 108
rect 79 70 113 111
rect -417 58 -351 70
rect -417 -58 -410 58
rect -358 -58 -351 58
rect -311 58 -265 70
rect -311 0 -305 58
rect -417 -70 -351 -58
rect -319 -9 -305 0
rect -271 0 -265 58
rect -225 61 -159 70
rect -225 9 -218 61
rect -166 9 -159 61
rect -225 0 -209 9
rect -271 -9 -257 0
rect -319 -61 -314 -9
rect -262 -61 -257 -9
rect -319 -70 -257 -61
rect -215 -58 -209 0
rect -175 0 -159 9
rect -119 58 -73 70
rect -119 0 -113 58
rect -175 -58 -169 0
rect -215 -70 -169 -58
rect -127 -9 -113 0
rect -79 0 -73 58
rect -33 58 33 70
rect -79 -9 -65 0
rect -127 -61 -122 -9
rect -70 -61 -65 -9
rect -127 -70 -65 -61
rect -33 -58 -26 58
rect 26 -58 33 58
rect 65 62 127 70
rect 65 10 70 62
rect 122 10 127 62
rect 65 0 79 10
rect -33 -70 33 -58
rect 73 -58 79 0
rect 113 0 127 10
rect 169 58 215 70
rect 169 0 175 58
rect 113 -58 119 0
rect 73 -70 119 -58
rect 159 -9 175 0
rect 209 0 215 58
rect 257 61 319 70
rect 257 9 262 61
rect 314 9 319 61
rect 257 0 271 9
rect 209 -9 225 0
rect 159 -61 166 -9
rect 218 -61 225 -9
rect 159 -70 225 -61
rect 265 -58 271 0
rect 305 0 319 9
rect 351 58 417 70
rect 305 -58 311 0
rect 265 -70 311 -58
rect 351 -58 358 58
rect 410 -58 417 58
rect 351 -70 417 -58
rect -113 -111 -79 -70
rect 310 -108 362 -102
rect -365 -117 -307 -111
rect -365 -151 -353 -117
rect -319 -151 -307 -117
rect -365 -157 -307 -151
rect -173 -117 -79 -111
rect 19 -117 77 -111
rect -173 -151 -161 -117
rect -127 -151 31 -117
rect 65 -151 77 -117
rect -173 -157 -115 -151
rect 19 -157 77 -151
rect 211 -117 269 -111
rect 211 -151 223 -117
rect 257 -151 310 -117
rect 211 -157 269 -151
rect 310 -166 362 -160
<< via1 >>
rect -362 108 -310 160
rect -410 -58 -401 58
rect -401 -58 -367 58
rect -367 -58 -358 58
rect -218 58 -166 61
rect -218 9 -209 58
rect -209 9 -175 58
rect -175 9 -166 58
rect -314 -58 -305 -9
rect -305 -58 -271 -9
rect -271 -58 -262 -9
rect -314 -61 -262 -58
rect -122 -58 -113 -9
rect -113 -58 -79 -9
rect -79 -58 -70 -9
rect -122 -61 -70 -58
rect -26 -58 -17 58
rect -17 -58 17 58
rect 17 -58 26 58
rect 70 58 122 62
rect 70 10 79 58
rect 79 10 113 58
rect 113 10 122 58
rect 262 58 314 61
rect 262 9 271 58
rect 271 9 305 58
rect 305 9 314 58
rect 166 -58 175 -9
rect 175 -58 209 -9
rect 209 -58 218 -9
rect 166 -61 218 -58
rect 358 -58 367 58
rect 367 -58 401 58
rect 401 -58 410 58
rect 310 -160 362 -108
<< metal2 >>
rect -551 151 -517 253
rect -368 151 -362 160
rect -551 117 -362 151
rect -368 108 -362 117
rect -310 108 -304 160
rect -417 58 -351 70
rect -417 -58 -412 58
rect -356 -58 -351 58
rect -229 63 -155 72
rect -229 7 -220 63
rect -164 7 -155 63
rect -417 -70 -351 -58
rect -319 -9 -257 0
rect -229 -2 -155 7
rect -33 58 33 70
rect -319 -61 -314 -9
rect -262 -36 -257 -9
rect -127 -9 -65 0
rect -127 -36 -122 -9
rect -262 -61 -122 -36
rect -70 -61 -65 -9
rect -319 -70 -65 -61
rect -33 -58 -28 58
rect 28 -58 33 58
rect 65 62 319 70
rect 65 10 70 62
rect 122 61 319 62
rect 122 36 262 61
rect 122 10 127 36
rect 65 0 127 10
rect 257 9 262 36
rect 314 9 319 61
rect -33 -70 33 -58
rect 155 -7 229 2
rect 257 0 319 9
rect 351 58 417 70
rect 155 -63 164 -7
rect 220 -63 229 -7
rect 155 -72 229 -63
rect 351 -58 356 58
rect 412 -58 417 58
rect 351 -70 417 -58
rect 304 -160 310 -108
rect 362 -117 368 -108
rect 517 -117 551 253
rect 362 -151 551 -117
rect 362 -160 368 -151
<< via2 >>
rect -412 -58 -410 58
rect -410 -58 -358 58
rect -358 -58 -356 58
rect -220 61 -164 63
rect -220 9 -218 61
rect -218 9 -166 61
rect -166 9 -164 61
rect -220 7 -164 9
rect -28 -58 -26 58
rect -26 -58 26 58
rect 26 -58 28 58
rect 164 -9 220 -7
rect 164 -61 166 -9
rect 166 -61 218 -9
rect 218 -61 220 -9
rect 164 -63 220 -61
rect 356 -58 358 58
rect 358 -58 410 58
rect 410 -58 412 58
<< metal3 >>
rect -417 63 33 72
rect -417 58 -220 63
rect -417 -58 -412 58
rect -356 12 -220 58
rect -356 -58 -351 12
rect -229 7 -220 12
rect -164 58 33 63
rect -164 12 -28 58
rect -164 7 -155 12
rect -229 -2 -155 7
rect -417 -70 -351 -58
rect -33 -58 -28 12
rect 28 -12 33 58
rect 351 58 417 72
rect 155 -7 229 2
rect 155 -12 164 -7
rect 28 -58 164 -12
rect -33 -63 164 -58
rect 220 -12 229 -7
rect 351 -12 356 58
rect 220 -58 356 -12
rect 412 -58 417 58
rect 220 -63 417 -58
rect -33 -70 417 -63
rect -414 -72 -351 -70
rect -30 -72 417 -70
<< properties >>
string FIXED_BBOX -498 -236 498 236
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.7 l 0.15 m 1 nf 8 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
