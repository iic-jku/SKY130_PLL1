magic
tech sky130A
magscale 1 2
timestamp 1668153059
<< pwell >>
rect -551 -280 551 280
<< nmos >>
rect -351 -70 -321 70
rect -255 -70 -225 70
rect -159 -70 -129 70
rect -63 -70 -33 70
rect 33 -70 63 70
rect 129 -70 159 70
rect 225 -70 255 70
rect 321 -70 351 70
<< ndiff >>
rect -413 58 -351 70
rect -413 -58 -401 58
rect -367 -58 -351 58
rect -413 -70 -351 -58
rect -321 58 -255 70
rect -321 -58 -305 58
rect -271 -58 -255 58
rect -321 -70 -255 -58
rect -225 58 -159 70
rect -225 -58 -209 58
rect -175 -58 -159 58
rect -225 -70 -159 -58
rect -129 58 -63 70
rect -129 -58 -113 58
rect -79 -58 -63 58
rect -129 -70 -63 -58
rect -33 58 33 70
rect -33 -58 -17 58
rect 17 -58 33 58
rect -33 -70 33 -58
rect 63 58 129 70
rect 63 -58 79 58
rect 113 -58 129 58
rect 63 -70 129 -58
rect 159 58 225 70
rect 159 -58 175 58
rect 209 -58 225 58
rect 159 -70 225 -58
rect 255 58 321 70
rect 255 -58 271 58
rect 305 -58 321 58
rect 255 -70 321 -58
rect 351 58 413 70
rect 351 -58 367 58
rect 401 -58 413 58
rect 351 -70 413 -58
<< ndiffc >>
rect -401 -58 -367 58
rect -305 -58 -271 58
rect -209 -58 -175 58
rect -113 -58 -79 58
rect -17 -58 17 58
rect 79 -58 113 58
rect 175 -58 209 58
rect 271 -58 305 58
rect 367 -58 401 58
<< psubdiff >>
rect -515 210 -419 244
rect 419 210 515 244
rect -515 148 -481 210
rect 481 148 515 210
rect -515 -210 -481 -148
rect 481 -210 515 -148
rect -515 -244 -419 -210
rect 419 -244 515 -210
<< psubdiffcont >>
rect -419 210 419 244
rect -515 -148 -481 148
rect 481 -148 515 148
rect -419 -244 419 -210
<< poly >>
rect -273 142 273 158
rect -273 108 -257 142
rect -223 108 -161 142
rect -127 108 -65 142
rect -31 108 31 142
rect 65 108 127 142
rect 161 108 223 142
rect 257 108 273 142
rect -351 70 -321 96
rect -273 92 273 108
rect -255 70 -225 92
rect -159 70 -129 92
rect -63 70 -33 92
rect 33 70 63 92
rect 129 70 159 92
rect 225 70 255 92
rect 321 70 351 96
rect -351 -92 -321 -70
rect -369 -108 -303 -92
rect -255 -96 -225 -70
rect -159 -96 -129 -70
rect -63 -96 -33 -70
rect 33 -96 63 -70
rect 129 -96 159 -70
rect 225 -96 255 -70
rect 321 -92 351 -70
rect -369 -142 -353 -108
rect -319 -142 -303 -108
rect -369 -158 -303 -142
rect 303 -108 369 -92
rect 303 -142 319 -108
rect 353 -142 369 -108
rect 303 -158 369 -142
<< polycont >>
rect -257 108 -223 142
rect -161 108 -127 142
rect -65 108 -31 142
rect 31 108 65 142
rect 127 108 161 142
rect 223 108 257 142
rect -353 -142 -319 -108
rect 319 -142 353 -108
<< locali >>
rect -515 210 -419 244
rect 419 210 515 244
rect -515 148 -481 210
rect 481 148 515 210
rect -273 108 -257 142
rect -223 108 -161 142
rect -127 108 -65 142
rect -31 108 31 142
rect 65 108 127 142
rect 161 108 223 142
rect 257 108 273 142
rect -515 -210 -481 -148
rect -401 58 -367 74
rect -401 -108 -367 -58
rect -305 58 -271 74
rect -305 -74 -271 -58
rect -209 58 -175 74
rect -209 -74 -175 -58
rect -113 58 -79 74
rect -113 -74 -79 -58
rect -17 58 17 74
rect -17 -74 17 -58
rect 79 58 113 74
rect 79 -74 113 -58
rect 175 58 209 74
rect 175 -74 209 -58
rect 271 58 305 74
rect 271 -74 305 -58
rect 367 58 401 74
rect 367 -108 401 -58
rect -401 -142 -353 -108
rect -319 -142 -303 -108
rect 303 -142 319 -108
rect 353 -142 401 -108
rect -401 -210 -367 -142
rect 367 -210 401 -142
rect 481 -210 515 -148
rect -515 -244 -419 -210
rect 419 -244 515 -210
<< viali >>
rect -257 108 -223 142
rect -161 108 -127 142
rect -65 108 -31 142
rect 31 108 65 142
rect 127 108 161 142
rect 223 108 257 142
rect -401 -58 -367 58
rect -305 -58 -271 58
rect -209 -58 -175 58
rect -113 -58 -79 58
rect -17 -58 17 58
rect 79 -58 113 58
rect 175 -58 209 58
rect 271 -58 305 58
rect 367 -58 401 58
rect -353 -142 -319 -108
rect 319 -142 353 -108
<< metal1 >>
rect -269 142 -211 148
rect -173 142 -115 148
rect -77 142 -19 148
rect 19 142 77 148
rect 115 142 173 148
rect 211 142 269 148
rect -273 108 -257 142
rect -223 108 -161 142
rect -127 108 -65 142
rect -31 108 31 142
rect 65 108 127 142
rect 161 108 223 142
rect 257 108 273 142
rect -269 102 -211 108
rect -173 102 -115 108
rect -77 102 -19 108
rect 19 102 77 108
rect 115 102 173 108
rect 211 102 269 108
rect -407 58 -361 70
rect -407 -1 -401 58
rect -413 -8 -401 -1
rect -367 -1 -361 58
rect -311 58 -265 70
rect -311 -1 -305 58
rect -367 -8 -305 -1
rect -271 -1 -265 58
rect -221 63 -163 70
rect -221 7 -219 63
rect -165 7 -163 63
rect -221 0 -209 7
rect -271 -8 -259 -1
rect -413 -64 -411 -8
rect -357 -64 -315 -8
rect -261 -64 -259 -8
rect -413 -70 -259 -64
rect -215 -58 -209 0
rect -175 0 -163 7
rect -119 58 -73 70
rect -175 -58 -169 0
rect -119 -1 -113 58
rect -215 -70 -169 -58
rect -125 -8 -113 -1
rect -79 -1 -73 58
rect -29 63 29 70
rect -29 7 -27 63
rect 27 7 29 63
rect -29 0 -17 7
rect -79 -8 -67 -1
rect -125 -64 -123 -8
rect -69 -64 -67 -8
rect -125 -70 -67 -64
rect -23 -58 -17 0
rect 17 0 29 7
rect 73 58 119 70
rect 17 -58 23 0
rect 73 -1 79 58
rect -23 -70 23 -58
rect 67 -8 79 -1
rect 113 -1 119 58
rect 163 63 221 70
rect 163 7 165 63
rect 219 7 221 63
rect 163 0 175 7
rect 113 -8 125 -1
rect 67 -64 69 -8
rect 123 -64 125 -8
rect 67 -70 125 -64
rect 169 -58 175 0
rect 209 0 221 7
rect 265 58 311 70
rect 209 -58 215 0
rect 265 -1 271 58
rect 169 -70 215 -58
rect 259 -8 271 -1
rect 305 -1 311 58
rect 361 58 407 70
rect 361 -1 367 58
rect 305 -8 367 -1
rect 401 -1 407 58
rect 401 -8 413 -1
rect 259 -64 261 -8
rect 315 -64 357 -8
rect 411 -64 413 -8
rect 259 -70 413 -64
rect -401 -102 -365 -70
rect 365 -102 401 -70
rect -401 -108 -307 -102
rect -401 -142 -353 -108
rect -319 -142 -307 -108
rect -401 -148 -307 -142
rect 307 -108 401 -102
rect 307 -142 319 -108
rect 353 -142 401 -108
rect 307 -148 401 -142
<< via1 >>
rect -219 58 -165 63
rect -219 7 -209 58
rect -209 7 -175 58
rect -175 7 -165 58
rect -411 -58 -401 -8
rect -401 -58 -367 -8
rect -367 -58 -357 -8
rect -411 -64 -357 -58
rect -315 -58 -305 -8
rect -305 -58 -271 -8
rect -271 -58 -261 -8
rect -315 -64 -261 -58
rect -27 58 27 63
rect -27 7 -17 58
rect -17 7 17 58
rect 17 7 27 58
rect -123 -58 -113 -8
rect -113 -58 -79 -8
rect -79 -58 -69 -8
rect -123 -64 -69 -58
rect 165 58 219 63
rect 165 7 175 58
rect 175 7 209 58
rect 209 7 219 58
rect 69 -58 79 -8
rect 79 -58 113 -8
rect 113 -58 123 -8
rect 69 -64 123 -58
rect 261 -58 271 -8
rect 271 -58 305 -8
rect 305 -58 315 -8
rect 261 -64 315 -58
rect 357 -58 367 -8
rect 367 -58 401 -8
rect 401 -58 411 -8
rect 357 -64 411 -58
<< metal2 >>
rect -221 63 225 70
rect -221 7 -219 63
rect -165 28 -27 63
rect -165 7 -163 28
rect -221 0 -163 7
rect -29 7 -27 28
rect 27 28 165 63
rect 27 7 29 28
rect -29 0 29 7
rect 163 7 165 28
rect 219 28 225 63
rect 219 7 221 28
rect 163 0 221 7
rect -413 -8 -259 -1
rect -413 -64 -411 -8
rect -357 -64 -315 -8
rect -261 -29 -259 -8
rect -125 -8 -67 -1
rect -125 -29 -123 -8
rect -261 -64 -123 -29
rect -69 -29 -67 -8
rect 67 -8 125 -1
rect 67 -29 69 -8
rect -69 -64 69 -29
rect 123 -29 125 -8
rect 259 -8 413 -1
rect 259 -29 261 -8
rect 123 -64 261 -29
rect 315 -64 357 -8
rect 411 -64 413 -8
rect -413 -70 413 -64
<< properties >>
string FIXED_BBOX -498 -227 498 227
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.7 l 0.150 m 1 nf 8 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
