magic
tech sky130A
magscale 1 2
timestamp 1659940462
<< error_p >>
rect -365 -108 -307 -102
rect 307 -108 365 -102
rect -365 -142 -353 -108
rect 307 -142 319 -108
rect -365 -148 -307 -142
rect 307 -148 365 -142
<< pwell >>
rect -551 -280 551 280
<< nmos >>
rect -351 -70 -321 70
rect -255 -70 -225 70
rect -159 -70 -129 70
rect -63 -70 -33 70
rect 33 -70 63 70
rect 129 -70 159 70
rect 225 -70 255 70
rect 321 -70 351 70
<< ndiff >>
rect -413 58 -351 70
rect -413 2 -401 58
rect -421 -58 -401 2
rect -367 -58 -351 58
rect -421 -70 -351 -58
rect -321 58 -255 70
rect -321 -58 -305 58
rect -271 -58 -255 58
rect -321 -70 -255 -58
rect -225 58 -159 70
rect -225 -58 -209 58
rect -175 -58 -159 58
rect -225 -70 -159 -58
rect -129 58 -63 70
rect -129 -58 -113 58
rect -79 -58 -63 58
rect -129 -70 -63 -58
rect -33 58 33 70
rect -33 -58 -17 58
rect 17 -58 33 58
rect -33 -70 33 -58
rect 63 58 129 70
rect 63 -58 79 58
rect 113 -58 129 58
rect 63 -70 129 -58
rect 159 58 225 70
rect 159 -58 175 58
rect 209 -58 225 58
rect 159 -70 225 -58
rect 255 58 321 70
rect 255 -58 271 58
rect 305 -58 321 58
rect 255 -70 321 -58
rect 351 58 413 70
rect 351 -58 367 58
rect 401 2 413 58
rect 401 -58 421 2
rect 351 -70 421 -58
<< ndiffc >>
rect -401 -58 -367 58
rect -305 -58 -271 58
rect -209 -58 -175 58
rect -113 -58 -79 58
rect -17 -58 17 58
rect 79 -58 113 58
rect 175 -58 209 58
rect 271 -58 305 58
rect 367 -58 401 58
<< psubdiff >>
rect -515 210 -419 244
rect 419 210 515 244
rect -515 148 -481 210
rect 481 148 515 210
rect -515 -210 -481 -148
rect 481 -210 515 -148
rect -515 -244 -419 -210
rect 419 -244 515 -210
<< psubdiffcont >>
rect -419 210 419 244
rect -515 -148 -481 148
rect 481 -148 515 148
rect -419 -244 419 -210
<< poly >>
rect -273 142 273 158
rect -273 108 -257 142
rect -223 108 -161 142
rect -127 108 -65 142
rect -31 108 31 142
rect 65 108 127 142
rect 161 108 223 142
rect 257 108 273 142
rect -351 70 -321 96
rect -273 92 273 108
rect -255 70 -225 92
rect -159 70 -129 92
rect -63 70 -33 92
rect 33 70 63 92
rect 129 70 159 92
rect 225 70 255 92
rect 321 70 351 96
rect -351 -92 -321 -70
rect -369 -108 -303 -92
rect -255 -96 -225 -70
rect -159 -96 -129 -70
rect -63 -96 -33 -70
rect 33 -96 63 -70
rect 129 -96 159 -70
rect 225 -96 255 -70
rect 321 -92 351 -70
rect -369 -142 -353 -108
rect -319 -142 -303 -108
rect -369 -158 -303 -142
rect 303 -108 369 -92
rect 303 -142 319 -108
rect 353 -142 369 -108
rect 303 -158 369 -142
<< polycont >>
rect -257 108 -223 142
rect -161 108 -127 142
rect -65 108 -31 142
rect 31 108 65 142
rect 127 108 161 142
rect 223 108 257 142
rect -353 -142 -319 -108
rect 319 -142 353 -108
<< locali >>
rect -515 210 -419 244
rect 419 210 515 244
rect -515 148 -481 210
rect 481 148 515 210
rect -273 108 -257 142
rect -223 108 -161 142
rect -127 108 -65 142
rect -31 108 31 142
rect 65 108 127 142
rect 161 108 223 142
rect 257 108 273 142
rect -401 58 -367 74
rect -401 -74 -367 -58
rect -305 58 -271 74
rect -305 -74 -271 -58
rect -209 58 -175 74
rect -209 -74 -175 -58
rect -113 58 -79 74
rect -113 -74 -79 -58
rect -17 58 17 74
rect -17 -74 17 -58
rect 79 58 113 74
rect 79 -74 113 -58
rect 175 58 209 74
rect 175 -74 209 -58
rect 271 58 305 74
rect 271 -74 305 -58
rect 367 58 401 74
rect 367 -74 401 -58
rect -369 -142 -353 -108
rect -319 -142 -303 -108
rect 303 -142 319 -108
rect 353 -142 369 -108
rect -515 -210 -481 -148
rect 551 -95 621 -25
rect 481 -210 515 -148
rect -515 -244 -419 -210
rect 419 -244 515 -210
<< viali >>
rect -257 108 -223 142
rect -161 108 -127 142
rect -65 108 -31 142
rect 31 108 65 142
rect 127 108 161 142
rect 223 108 257 142
rect -401 -58 -367 58
rect -305 -58 -271 58
rect -209 -58 -175 58
rect -113 -58 -79 58
rect -17 -58 17 58
rect 79 -58 113 58
rect 175 -58 209 58
rect 271 -58 305 58
rect 367 -58 401 58
rect -353 -142 -319 -108
rect 319 -142 353 -108
<< metal1 >>
rect -269 142 -211 148
rect -173 142 -115 148
rect -77 142 -19 148
rect 19 142 77 148
rect 115 142 173 148
rect 211 142 269 148
rect -269 108 -257 142
rect -223 108 -161 142
rect -127 108 -65 142
rect -31 108 31 142
rect 65 108 127 142
rect 161 108 223 142
rect 257 108 269 142
rect -269 102 -211 108
rect -173 102 -115 108
rect -77 102 -19 108
rect 19 102 77 108
rect 115 102 173 108
rect 211 102 269 108
rect -407 58 -361 70
rect -407 0 -401 58
rect -414 -9 -401 0
rect -367 0 -361 58
rect -311 58 -265 70
rect -311 0 -305 58
rect -367 -9 -354 0
rect -414 -61 -410 -9
rect -358 -61 -354 -9
rect -414 -70 -354 -61
rect -318 -9 -305 0
rect -271 0 -265 58
rect -222 61 -162 70
rect -222 9 -218 61
rect -166 9 -162 61
rect -222 0 -209 9
rect -271 -9 -258 0
rect -318 -61 -314 -9
rect -262 -61 -258 -9
rect -318 -70 -258 -61
rect -215 -58 -209 0
rect -175 0 -162 9
rect -119 58 -73 70
rect -119 0 -113 58
rect -175 -58 -169 0
rect -215 -70 -169 -58
rect -126 -9 -113 0
rect -79 0 -73 58
rect -30 61 30 70
rect -30 9 -26 61
rect 26 9 30 61
rect -30 0 -17 9
rect -79 -9 -66 0
rect -126 -61 -122 -9
rect -70 -61 -66 -9
rect -126 -70 -66 -61
rect -23 -58 -17 0
rect 17 0 30 9
rect 73 58 119 70
rect 73 0 79 58
rect 17 -58 23 0
rect -23 -70 23 -58
rect 66 -9 79 0
rect 113 0 119 58
rect 162 61 222 70
rect 162 9 166 61
rect 218 9 222 61
rect 162 0 175 9
rect 113 -9 126 0
rect 66 -61 70 -9
rect 122 -61 126 -9
rect 66 -70 126 -61
rect 169 -58 175 0
rect 209 0 222 9
rect 265 58 311 70
rect 265 0 271 58
rect 209 -58 215 0
rect 169 -70 215 -58
rect 258 -9 271 0
rect 305 0 311 58
rect 361 58 407 70
rect 361 0 367 58
rect 305 -9 318 0
rect 258 -61 262 -9
rect 314 -61 318 -9
rect 258 -70 318 -61
rect 354 -9 367 0
rect 401 0 407 58
rect 401 -9 414 0
rect 354 -61 358 -9
rect 410 -61 414 -9
rect 354 -70 414 -61
rect -365 -108 -307 -102
rect -365 -142 -353 -108
rect -319 -142 -307 -108
rect -365 -148 -307 -142
rect 307 -108 365 -102
rect 307 -142 319 -108
rect 353 -142 365 -108
rect 307 -148 365 -142
<< via1 >>
rect -410 -58 -401 -9
rect -401 -58 -367 -9
rect -367 -58 -358 -9
rect -410 -61 -358 -58
rect -218 58 -166 61
rect -218 9 -209 58
rect -209 9 -175 58
rect -175 9 -166 58
rect -314 -58 -305 -9
rect -305 -58 -271 -9
rect -271 -58 -262 -9
rect -314 -61 -262 -58
rect -26 58 26 61
rect -26 9 -17 58
rect -17 9 17 58
rect 17 9 26 58
rect -122 -58 -113 -9
rect -113 -58 -79 -9
rect -79 -58 -70 -9
rect -122 -61 -70 -58
rect 166 58 218 61
rect 166 9 175 58
rect 175 9 209 58
rect 209 9 218 58
rect 70 -58 79 -9
rect 79 -58 113 -9
rect 113 -58 122 -9
rect 70 -61 122 -58
rect 262 -58 271 -9
rect 271 -58 305 -9
rect 305 -58 314 -9
rect 262 -61 314 -58
rect 358 -58 367 -9
rect 367 -58 401 -9
rect 401 -58 410 -9
rect 358 -61 410 -58
<< metal2 >>
rect -222 61 222 70
rect -222 9 -218 61
rect -166 36 -26 61
rect -166 9 -162 36
rect -421 -7 -251 2
rect -222 0 -162 9
rect -30 9 -26 36
rect 26 36 166 61
rect 26 9 30 36
rect -421 -63 -412 -7
rect -356 -63 -316 -7
rect -260 -63 -251 -7
rect -421 -72 -251 -63
rect -133 -7 -59 2
rect -30 0 30 9
rect 162 9 166 36
rect 218 9 222 61
rect -133 -63 -124 -7
rect -68 -63 -59 -7
rect -133 -72 -59 -63
rect 59 -7 133 2
rect 162 0 222 9
rect 59 -63 68 -7
rect 124 -63 133 -7
rect 59 -72 133 -63
rect 251 -7 421 2
rect 251 -63 260 -7
rect 316 -63 356 -7
rect 412 -63 421 -7
rect 251 -72 421 -63
<< via2 >>
rect -412 -9 -356 -7
rect -412 -61 -410 -9
rect -410 -61 -358 -9
rect -358 -61 -356 -9
rect -412 -63 -356 -61
rect -316 -9 -260 -7
rect -316 -61 -314 -9
rect -314 -61 -262 -9
rect -262 -61 -260 -9
rect -316 -63 -260 -61
rect -124 -9 -68 -7
rect -124 -61 -122 -9
rect -122 -61 -70 -9
rect -70 -61 -68 -9
rect -124 -63 -68 -61
rect 68 -9 124 -7
rect 68 -61 70 -9
rect 70 -61 122 -9
rect 122 -61 124 -9
rect 68 -63 124 -61
rect 260 -9 316 -7
rect 260 -61 262 -9
rect 262 -61 314 -9
rect 314 -61 316 -9
rect 260 -63 316 -61
rect 356 -9 412 -7
rect 356 -61 358 -9
rect 358 -61 410 -9
rect 410 -61 412 -9
rect 356 -63 412 -61
<< metal3 >>
rect -421 -7 -251 2
rect -421 -63 -412 -7
rect -356 -63 -316 -7
rect -260 -10 -251 -7
rect -133 -7 -59 2
rect -133 -10 -124 -7
rect -260 -63 -124 -10
rect -68 -10 -59 -7
rect 59 -7 133 2
rect 59 -10 68 -7
rect -68 -63 68 -10
rect 124 -10 133 -7
rect 251 -7 421 2
rect 251 -10 260 -7
rect 124 -63 260 -10
rect 316 -63 356 -7
rect 412 -63 421 -7
rect -421 -70 421 -63
rect -421 -72 -251 -70
rect -133 -72 -59 -70
rect 59 -72 133 -70
rect 251 -72 421 -70
<< properties >>
string FIXED_BBOX -498 -227 498 227
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.7 l 0.150 m 1 nf 8 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
