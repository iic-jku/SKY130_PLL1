magic
tech sky130A
magscale 1 2
timestamp 1665586327
<< metal1 >>
rect 7475 9287 8045 10023
rect 931 9269 1501 9287
rect 931 8872 947 9269
rect 1485 8872 1501 9269
rect 931 8855 1501 8872
rect 1749 9269 3137 9287
rect 1749 8872 2583 9269
rect 3121 8872 3137 9269
rect 1749 8855 3137 8872
rect 3385 9269 4773 9287
rect 3385 8872 4219 9269
rect 4757 8872 4773 9269
rect 3385 8855 4773 8872
rect 5021 9269 6409 9287
rect 5021 8872 5855 9269
rect 6393 8872 6409 9269
rect 5021 8855 6409 8872
rect 6657 8855 8045 9287
rect 931 4117 1501 5313
rect 1749 5296 2319 5313
rect 1749 4899 1765 5296
rect 2303 4899 2319 5296
rect 1749 4117 2319 4899
rect 2567 4117 3137 5313
rect 3385 4531 3955 4549
rect 3385 4134 3401 4531
rect 3939 4134 3955 4531
rect 3385 4117 3955 4134
rect 4203 4117 4773 5313
rect 5839 4117 6409 5313
rect 7475 4117 8045 5313
rect 1749 558 2319 575
rect 931 -593 1501 167
rect 1749 161 1765 558
rect 2303 161 2319 558
rect 3385 558 3955 575
rect 1749 143 2319 161
rect 2567 -593 3137 179
rect 3385 161 3401 558
rect 3939 161 3955 558
rect 3385 143 3955 161
rect 4203 -593 4773 167
rect 5839 -593 6409 176
rect 7475 -593 8045 176
<< via1 >>
rect 947 8872 1485 9269
rect 2583 8872 3121 9269
rect 4219 8872 4757 9269
rect 5855 8872 6393 9269
rect 1765 4899 2303 5296
rect 3401 4899 3939 5296
rect 3401 4134 3939 4531
rect 5037 4899 5575 5296
rect 6673 4899 7211 5296
rect 1765 161 2303 558
rect 3401 161 3939 558
<< metal2 >>
rect 931 9269 1501 9287
rect 931 8872 947 9269
rect 1485 8872 1501 9269
rect 931 5313 1501 8872
rect 2567 9269 3137 9287
rect 2567 8872 2583 9269
rect 3121 8872 3137 9269
rect 2567 5313 3137 8872
rect 4203 9269 4773 9287
rect 4203 8872 4219 9269
rect 4757 8872 4773 9269
rect 4203 5313 4773 8872
rect 5839 9269 6409 9287
rect 5839 8872 5855 9269
rect 6393 8872 6409 9269
rect 5839 5313 6409 8872
rect 931 5296 2319 5313
rect 931 4899 1765 5296
rect 2303 4899 2319 5296
rect 931 4881 2319 4899
rect 2567 5296 3955 5313
rect 2567 4899 3401 5296
rect 3939 4899 3955 5296
rect 2567 4881 3955 4899
rect 4203 5296 5591 5313
rect 4203 4899 5037 5296
rect 5575 4899 5591 5296
rect 4203 4881 5591 4899
rect 5839 5296 7227 5313
rect 5839 4899 6673 5296
rect 7211 4899 7227 5296
rect 5839 4881 7227 4899
rect -485 4531 3955 4549
rect -485 4134 3401 4531
rect 3939 4134 3955 4531
rect -485 4117 3955 4134
rect 1749 558 3955 575
rect 1749 161 1765 558
rect 2303 161 3401 558
rect 3939 161 3955 558
rect 1749 143 3955 161
use sky130_fd_pr__res_high_po_2p85_DZG53T  sky130_fd_pr__res_high_po_2p85_DZG53T_0
timestamp 1665586327
transform 1 0 4488 0 1 7084
box -4541 -2369 4541 2369
use sky130_fd_pr__res_high_po_2p85_DZG53T  sky130_fd_pr__res_high_po_2p85_DZG53T_1
timestamp 1665586327
transform 1 0 4488 0 1 2346
box -4541 -2369 4541 2369
<< labels >>
rlabel metal1 931 -593 1501 -23 3 b0
rlabel metal1 2567 -593 3137 -23 3 b1
rlabel metal1 4203 -593 4773 -23 0 b2
rlabel metal1 5839 -593 6409 -23 5 b3
rlabel metal1 7475 -593 8045 -23 0 b4
rlabel metal2 -485 4117 -53 4549 7 vss
rlabel metal1 7475 9453 8045 10023 0 vout
<< end >>
