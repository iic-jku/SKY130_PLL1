magic
tech sky130A
magscale 1 2
timestamp 1668332298
<< nwell >>
rect 1530 -5003 1739 -4682
rect 3804 -5003 4125 -4682
rect 6301 -5003 6511 -4680
rect 1209 -6934 1765 -6613
rect 3594 -6934 4478 -6613
rect 5966 -6932 6832 -6611
<< metal1 >>
rect 2170 6916 2212 6976
rect 3290 6917 3332 6976
rect 4704 6917 4746 6976
rect 2150 6901 2232 6916
rect 2150 6849 2165 6901
rect 2217 6849 2232 6901
rect 2150 6834 2232 6849
rect 3270 6901 3352 6917
rect 3270 6849 3285 6901
rect 3337 6849 3352 6901
rect 3270 6834 3352 6849
rect 4684 6901 4766 6917
rect 5824 6916 5866 6976
rect 4684 6849 4699 6901
rect 4751 6849 4766 6901
rect 4684 6834 4766 6849
rect 5804 6901 5886 6916
rect 5804 6849 5819 6901
rect 5871 6849 5886 6901
rect 5804 6834 5886 6849
rect 3597 6777 3677 6786
rect 3597 6595 3608 6777
rect 3660 6595 3677 6777
rect 3597 6586 3677 6595
rect 4352 6777 4458 6786
rect 4352 6595 4374 6777
rect 4426 6595 4458 6777
rect 4352 6586 4458 6595
rect 6120 6777 6226 6786
rect 6120 6595 6142 6777
rect 6194 6595 6226 6777
rect 6120 6586 6226 6595
rect 379 6416 579 6422
rect -755 6403 -703 6409
rect -755 6345 -703 6351
rect -750 6188 -708 6345
rect 2468 6407 2548 6416
rect 2468 6225 2479 6407
rect 2531 6225 2548 6407
rect 2468 6216 2548 6225
rect 2958 6407 3038 6416
rect 2958 6225 2969 6407
rect 3021 6225 3038 6407
rect 2958 6216 3038 6225
rect 4991 6407 5097 6416
rect 4991 6225 5013 6407
rect 5065 6225 5097 6407
rect 4991 6216 5097 6225
rect 5481 6407 5587 6416
rect 5481 6225 5503 6407
rect 5555 6225 5587 6407
rect 5481 6216 5587 6225
rect 7658 6216 7664 6416
rect 8740 6407 8792 6413
rect 8740 6349 8792 6355
rect 379 6210 579 6216
rect 8745 6177 8787 6349
rect 9 6154 209 6162
rect 9 6102 18 6154
rect 200 6102 209 6154
rect 9 6092 209 6102
rect 7828 6143 8028 6151
rect 7828 6091 7837 6143
rect 8019 6091 8028 6143
rect 7828 6081 8028 6091
rect 9 4155 209 4163
rect 9 4103 18 4155
rect 200 4103 209 4155
rect 9 4093 209 4103
rect 7828 4147 8028 4155
rect 7828 4095 7837 4147
rect 8019 4095 8028 4147
rect 7828 4085 8028 4095
rect 379 3909 579 3917
rect 379 3857 388 3909
rect 570 3857 579 3909
rect 379 3847 579 3857
rect 7458 3916 7658 3924
rect 7458 3864 7467 3916
rect 7649 3864 7658 3916
rect 7458 3854 7658 3864
rect 4122 3496 4128 3548
rect 4180 3496 4186 3548
rect 3986 3237 3992 3289
rect 4044 3237 4050 3289
rect 3850 3106 3856 3158
rect 3908 3106 3914 3158
rect 9 2632 209 2832
rect 379 2629 579 2829
rect 10780 771 10822 813
rect 2471 561 2541 570
rect 2471 379 2479 561
rect 2531 379 2541 561
rect 2471 370 2541 379
rect 2961 561 3031 570
rect 2961 379 2969 561
rect 3021 379 3031 561
rect 2961 370 3031 379
rect 5005 561 5075 570
rect 5005 379 5013 561
rect 5065 379 5075 561
rect 5005 370 5075 379
rect 5495 561 5565 570
rect 5495 379 5503 561
rect 5555 379 5565 561
rect 5495 370 5565 379
rect 7452 370 7458 570
rect 7658 370 7664 570
rect 1818 191 1929 200
rect 1818 9 1840 191
rect 1892 9 1929 191
rect 1818 0 1929 9
rect 3600 191 3670 200
rect 3600 9 3608 191
rect 3660 9 3670 191
rect 3600 0 3670 9
rect 4366 191 4436 200
rect 4366 9 4374 191
rect 4426 9 4436 191
rect 4366 0 4436 9
rect 6134 191 6204 200
rect 6134 9 6142 191
rect 6194 9 6204 191
rect 6134 0 6204 9
rect 2150 -63 2232 -48
rect 2150 -115 2165 -63
rect 2217 -115 2232 -63
rect 2150 -130 2232 -115
rect 3270 -63 3352 -48
rect 3270 -115 3285 -63
rect 3337 -115 3352 -63
rect 2170 -190 2212 -130
rect 3270 -131 3352 -115
rect 4684 -63 4766 -48
rect 4684 -115 4699 -63
rect 4751 -115 4766 -63
rect 4684 -131 4766 -115
rect 5804 -63 5886 -48
rect 5804 -115 5819 -63
rect 5871 -115 5886 -63
rect 5804 -130 5886 -115
rect 3290 -190 3332 -131
rect 4704 -190 4746 -131
rect 5824 -190 5866 -130
rect 7828 -303 8028 200
rect 7828 -362 7834 -303
rect 8021 -362 8028 -303
rect 7828 -367 8028 -362
rect 2170 -1027 2212 -1016
rect 5824 -1025 5866 -1016
rect 2165 -1033 2217 -1027
rect 2165 -1091 2217 -1085
rect 5819 -1031 5871 -1025
rect 5819 -1089 5871 -1083
rect 2170 -1100 2212 -1091
rect 5824 -1100 5866 -1089
rect 1492 -4768 1777 -4671
rect 3877 -4768 4163 -4671
rect 6262 -4766 6549 -4670
rect 3876 -5216 4162 -5215
rect 3876 -5312 4163 -5216
rect 1492 -6400 1777 -6303
rect 3877 -6400 4164 -6304
rect 6262 -6399 6549 -6303
rect 1492 -6944 1777 -6847
rect 3877 -6944 4164 -6848
rect 6263 -6943 6550 -6847
rect 1178 -7139 1530 -7099
rect 3564 -7139 3915 -7099
rect 4125 -7139 4476 -7099
rect 6511 -7137 6862 -7097
rect 1140 -7488 1777 -7392
rect 3525 -7488 4516 -7392
rect 6263 -7488 6902 -7392
<< via1 >>
rect 2165 6849 2217 6901
rect 3285 6849 3337 6901
rect 4699 6849 4751 6901
rect 5819 6849 5871 6901
rect 1840 6595 1892 6777
rect 3608 6595 3660 6777
rect 4374 6595 4426 6777
rect 6142 6595 6194 6777
rect -755 6351 -703 6403
rect 379 6216 579 6416
rect 2479 6225 2531 6407
rect 2969 6225 3021 6407
rect 5013 6225 5065 6407
rect 5503 6225 5555 6407
rect 7458 6216 7658 6416
rect 8740 6355 8792 6407
rect 18 6102 200 6154
rect 7837 6091 8019 6143
rect 18 4103 200 4155
rect 7837 4095 8019 4147
rect 388 3857 570 3909
rect 7467 3864 7649 3916
rect 4128 3496 4180 3548
rect 3992 3237 4044 3289
rect 3856 3106 3908 3158
rect 2479 379 2531 561
rect 2969 379 3021 561
rect 5013 379 5065 561
rect 5503 379 5555 561
rect 7458 370 7658 570
rect 1840 9 1892 191
rect 3608 9 3660 191
rect 4374 9 4426 191
rect 6142 9 6194 191
rect 2165 -115 2217 -63
rect 3285 -115 3337 -63
rect 4699 -115 4751 -63
rect 5819 -115 5871 -63
rect 7834 -362 8021 -303
rect 2165 -1085 2217 -1033
rect 5819 -1083 5871 -1031
<< metal2 >>
rect -750 8383 2212 8425
rect -750 6403 -708 8383
rect 2170 7844 2212 8383
rect 4704 7906 8787 7948
rect 4704 7802 4746 7906
rect 1832 6777 1902 7073
rect 2150 6905 2232 6916
rect 2150 6845 2161 6905
rect 2221 6845 2232 6905
rect 2150 6834 2232 6845
rect 1832 6595 1840 6777
rect 1892 6595 1902 6777
rect 1832 6586 1902 6595
rect 379 6416 579 6426
rect -761 6351 -755 6403
rect -703 6351 -697 6403
rect 373 6300 379 6416
rect -1079 6230 379 6300
rect -1079 5996 -1009 6230
rect 373 6216 379 6230
rect 579 6216 585 6416
rect 2471 6407 2541 7168
rect 2471 6225 2479 6407
rect 2531 6225 2541 6407
rect 2471 6216 2541 6225
rect 2961 6407 3031 7168
rect 3270 6905 3352 6917
rect 3270 6845 3281 6905
rect 3341 6845 3352 6905
rect 3270 6834 3352 6845
rect 3600 6777 3670 7072
rect 3600 6595 3608 6777
rect 3660 6595 3670 6777
rect 3600 6586 3670 6595
rect 4366 6777 4436 7072
rect 4684 6905 4766 6917
rect 4684 6845 4695 6905
rect 4755 6845 4766 6905
rect 4684 6834 4766 6845
rect 4366 6595 4374 6777
rect 4426 6595 4436 6777
rect 4366 6586 4436 6595
rect 2961 6225 2969 6407
rect 3021 6225 3031 6407
rect 2961 6216 3031 6225
rect 5005 6407 5075 7168
rect 5005 6225 5013 6407
rect 5065 6225 5075 6407
rect 5005 6216 5075 6225
rect 5495 6407 5565 7168
rect 5804 6905 5886 6916
rect 5804 6845 5815 6905
rect 5875 6845 5886 6905
rect 5804 6834 5886 6845
rect 6134 6777 6204 7072
rect 6134 6595 6142 6777
rect 6194 6595 6204 6777
rect 6134 6586 6204 6595
rect 5495 6225 5503 6407
rect 5555 6225 5565 6407
rect 5495 6216 5565 6225
rect 7458 6416 7658 6423
rect 8745 6407 8787 7906
rect 8734 6355 8740 6407
rect 8792 6355 8798 6407
rect 7658 6219 9116 6289
rect 7458 6210 7658 6216
rect -440 6154 209 6162
rect -440 6102 18 6154
rect 200 6102 209 6154
rect -440 6092 209 6102
rect 7828 6143 8477 6151
rect 7828 6091 7837 6143
rect 8019 6091 8477 6143
rect 7828 6081 8477 6091
rect 9046 5985 9116 6219
rect 9509 5294 9642 5328
rect -1079 3917 -1009 4355
rect -440 4155 209 4163
rect -440 4103 18 4155
rect 200 4103 209 4155
rect -440 4093 209 4103
rect 7828 4147 8477 4155
rect 7828 4095 7837 4147
rect 8019 4095 8477 4147
rect 7828 4085 8477 4095
rect 8407 4082 8477 4085
rect -750 4026 -708 4068
rect 8745 4030 8787 4057
rect -759 4017 -699 4026
rect -759 3948 -699 3957
rect 8736 4021 8796 4030
rect 8736 3952 8796 3961
rect 9046 3924 9116 4344
rect -1079 3909 579 3917
rect -1079 3857 388 3909
rect 570 3857 579 3909
rect -1079 3847 579 3857
rect 7458 3916 9116 3924
rect 7458 3864 7467 3916
rect 7649 3864 9116 3916
rect 7458 3854 9116 3864
rect 4128 3548 4180 3554
rect 9509 3539 9543 5294
rect 10562 5286 10864 5328
rect 4180 3505 9543 3539
rect 4128 3490 4180 3496
rect -1329 3363 2712 3423
rect 3979 3363 3988 3423
rect 4048 3363 4057 3423
rect 3992 3289 4044 3295
rect 4044 3246 9642 3280
rect 10561 3240 10864 3282
rect 3992 3231 4044 3237
rect 3856 3158 3908 3164
rect 3908 3115 9543 3149
rect 3856 3100 3908 3106
rect 9509 1232 9543 3115
rect 9509 1198 9642 1232
rect 10561 1194 10864 1236
rect 7458 570 7658 576
rect 2471 561 2541 570
rect 2471 379 2479 561
rect 2531 379 2541 561
rect 1832 191 1902 200
rect 1832 9 1840 191
rect 1892 9 1902 191
rect 1832 -286 1902 9
rect 2150 -59 2232 -48
rect 2150 -119 2161 -59
rect 2221 -119 2232 -59
rect 2150 -130 2232 -119
rect 2471 -382 2541 379
rect 2961 561 3031 570
rect 2961 379 2969 561
rect 3021 379 3031 561
rect 2961 -382 3031 379
rect 5005 561 5075 570
rect 5005 379 5013 561
rect 5065 379 5075 561
rect 3600 191 3670 200
rect 3600 9 3608 191
rect 3660 9 3670 191
rect 3270 -59 3352 -48
rect 3270 -119 3281 -59
rect 3341 -119 3352 -59
rect 3270 -131 3352 -119
rect 3600 -286 3670 9
rect 4366 191 4436 200
rect 4366 9 4374 191
rect 4426 9 4436 191
rect 4366 -286 4436 9
rect 4684 -59 4766 -48
rect 4684 -119 4695 -59
rect 4755 -119 4766 -59
rect 4684 -131 4766 -119
rect 5005 -382 5075 379
rect 5495 561 5565 570
rect 5495 379 5503 561
rect 5555 379 5565 561
rect 5495 -382 5565 379
rect 7658 370 7665 570
rect 7458 364 7658 370
rect 6134 191 6204 200
rect 6134 9 6142 191
rect 6194 9 6204 191
rect 5804 -59 5886 -48
rect 5804 -119 5815 -59
rect 5875 -119 5886 -59
rect 5804 -130 5886 -119
rect 6134 -286 6204 9
rect 7521 -21 7591 364
rect 7521 -91 9922 -21
rect 10491 -297 10561 -118
rect 7828 -303 10561 -297
rect 7828 -362 7834 -303
rect 8021 -362 10561 -303
rect 7828 -367 10561 -362
rect 1832 -1196 1902 -919
rect 2159 -1085 2165 -1033
rect 2217 -1085 2223 -1033
rect 2472 -1292 2541 -823
rect 5495 -1292 5564 -823
rect 5813 -1083 5819 -1031
rect 5871 -1083 5877 -1031
rect 6134 -1197 6204 -916
rect 2170 -3268 2212 -3220
rect 1696 -3333 2212 -3268
rect 5824 -3268 5866 -3220
rect 5824 -3333 6344 -3268
rect -771 -5071 -762 -5005
rect -696 -5071 -624 -5005
rect 1696 -5071 1761 -3333
rect 6279 -5071 6344 -3333
rect 8665 -5069 8733 -5003
rect 8799 -5069 8808 -5003
<< via2 >>
rect 2161 6901 2221 6905
rect 2161 6849 2165 6901
rect 2165 6849 2217 6901
rect 2217 6849 2221 6901
rect 2161 6845 2221 6849
rect 3281 6901 3341 6905
rect 3281 6849 3285 6901
rect 3285 6849 3337 6901
rect 3337 6849 3341 6901
rect 3281 6845 3341 6849
rect 4695 6901 4755 6905
rect 4695 6849 4699 6901
rect 4699 6849 4751 6901
rect 4751 6849 4755 6901
rect 4695 6845 4755 6849
rect 5815 6901 5875 6905
rect 5815 6849 5819 6901
rect 5819 6849 5871 6901
rect 5871 6849 5875 6901
rect 5815 6845 5875 6849
rect -759 3957 -699 4017
rect 8736 3961 8796 4021
rect 3988 3363 4048 3423
rect 2161 -63 2221 -59
rect 2161 -115 2165 -63
rect 2165 -115 2217 -63
rect 2217 -115 2221 -63
rect 2161 -119 2221 -115
rect 3281 -63 3341 -59
rect 3281 -115 3285 -63
rect 3285 -115 3337 -63
rect 3337 -115 3341 -63
rect 3281 -119 3341 -115
rect 4695 -63 4755 -59
rect 4695 -115 4699 -63
rect 4699 -115 4751 -63
rect 4751 -115 4755 -63
rect 4695 -119 4755 -115
rect 5815 -63 5875 -59
rect 5815 -115 5819 -63
rect 5819 -115 5871 -63
rect 5871 -115 5875 -63
rect 5815 -119 5875 -115
rect -762 -5071 -696 -5005
rect 8733 -5069 8799 -5003
<< metal3 >>
rect 2150 6910 2232 6916
rect 2150 6840 2156 6910
rect 2226 6840 2232 6910
rect 2150 6834 2232 6840
rect 3270 6910 3352 6917
rect 3270 6840 3276 6910
rect 3346 6840 3352 6910
rect 3270 6834 3352 6840
rect 4684 6910 4766 6917
rect 4684 6840 4690 6910
rect 4760 6840 4766 6910
rect 4684 6834 4766 6840
rect 5804 6910 5886 6916
rect 5804 6840 5810 6910
rect 5880 6840 5886 6910
rect 5804 6834 5886 6840
rect 2170 6786 2230 6834
rect 3272 6786 3332 6834
rect 4704 6786 4764 6834
rect 5806 6786 5866 6834
rect -764 4017 -694 4022
rect -764 3957 -759 4017
rect -699 3957 -694 4017
rect -764 3952 -694 3957
rect 8731 4021 8801 4026
rect 8731 3961 8736 4021
rect 8796 3961 8801 4021
rect 8731 3956 8801 3961
rect -759 -5000 -699 3952
rect 3983 3423 4053 3428
rect 3983 3363 3988 3423
rect 4048 3363 4053 3423
rect 3983 3358 4053 3363
rect 2170 -48 2230 0
rect 3272 -48 3332 0
rect 4704 -48 4764 0
rect 5806 -48 5866 0
rect 2150 -54 2232 -48
rect 2150 -124 2156 -54
rect 2226 -124 2232 -54
rect 2150 -130 2232 -124
rect 3270 -54 3352 -48
rect 3270 -124 3276 -54
rect 3346 -124 3352 -54
rect 3270 -131 3352 -124
rect 4684 -54 4766 -48
rect 4684 -124 4690 -54
rect 4760 -124 4766 -54
rect 4684 -131 4766 -124
rect 5804 -54 5886 -48
rect 5804 -124 5810 -54
rect 5880 -124 5886 -54
rect 5804 -130 5886 -124
rect 8736 -4998 8796 3956
rect -767 -5005 -691 -5000
rect -767 -5071 -762 -5005
rect -696 -5071 -691 -5005
rect -767 -5076 -691 -5071
rect 8728 -5003 8804 -4998
rect 8728 -5069 8733 -5003
rect 8799 -5069 8804 -5003
rect 8728 -5074 8804 -5069
<< via3 >>
rect 2156 6905 2226 6910
rect 2156 6845 2161 6905
rect 2161 6845 2221 6905
rect 2221 6845 2226 6905
rect 2156 6840 2226 6845
rect 3276 6905 3346 6910
rect 3276 6845 3281 6905
rect 3281 6845 3341 6905
rect 3341 6845 3346 6905
rect 3276 6840 3346 6845
rect 4690 6905 4760 6910
rect 4690 6845 4695 6905
rect 4695 6845 4755 6905
rect 4755 6845 4760 6905
rect 4690 6840 4760 6845
rect 5810 6905 5880 6910
rect 5810 6845 5815 6905
rect 5815 6845 5875 6905
rect 5875 6845 5880 6905
rect 5810 6840 5880 6845
rect 2156 -59 2226 -54
rect 2156 -119 2161 -59
rect 2161 -119 2221 -59
rect 2221 -119 2226 -59
rect 2156 -124 2226 -119
rect 3276 -59 3346 -54
rect 3276 -119 3281 -59
rect 3281 -119 3341 -59
rect 3341 -119 3346 -59
rect 3276 -124 3346 -119
rect 4690 -59 4760 -54
rect 4690 -119 4695 -59
rect 4695 -119 4755 -59
rect 4755 -119 4760 -59
rect 4690 -124 4760 -119
rect 5810 -59 5880 -54
rect 5810 -119 5815 -59
rect 5815 -119 5875 -59
rect 5875 -119 5880 -59
rect 5810 -124 5880 -119
<< metal4 >>
rect 2150 6910 2232 6916
rect 2150 6840 2156 6910
rect 2226 6840 2232 6910
rect 2150 6834 2232 6840
rect 3270 6910 3352 6917
rect 3270 6840 3276 6910
rect 3346 6840 3352 6910
rect 3270 6834 3352 6840
rect 4684 6910 4766 6917
rect 4684 6840 4690 6910
rect 4760 6840 4766 6910
rect 4684 6834 4766 6840
rect 5804 6910 5886 6916
rect 5804 6840 5810 6910
rect 5880 6840 5886 6910
rect 5804 6834 5886 6840
rect 2170 5703 2230 6834
rect 3272 5703 3332 6834
rect 4704 5702 4764 6834
rect 5806 5703 5866 6834
rect 2170 -48 2230 1083
rect 3272 -48 3332 1086
rect 4704 -48 4764 1083
rect 5806 -48 5866 1083
rect 2150 -54 2232 -48
rect 2150 -124 2156 -54
rect 2226 -124 2232 -54
rect 2150 -130 2232 -124
rect 3270 -54 3352 -48
rect 3270 -124 3276 -54
rect 3346 -124 3352 -54
rect 3270 -131 3352 -124
rect 4684 -54 4766 -48
rect 4684 -124 4690 -54
rect 4760 -124 4766 -54
rect 4684 -131 4766 -124
rect 5804 -54 5886 -48
rect 5804 -124 5810 -54
rect 5880 -124 5886 -54
rect 5804 -130 5886 -124
use d_ff_15  d_ff_15_0
timestamp 1668240031
transform -1 0 6263 0 1 -5264
box -98 -2224 2138 697
use d_ff_15  d_ff_15_1
timestamp 1668240031
transform -1 0 8649 0 1 -5262
box -98 -2224 2138 697
use d_ff_15  d_ff_15_2
timestamp 1668240031
transform 1 0 1777 0 1 -5264
box -98 -2224 2138 697
use d_ff_15  d_ff_15_3
timestamp 1668240031
transform 1 0 -608 0 1 -5264
box -98 -2224 2138 697
use inv_buffer2  inv_buffer2_0
timestamp 1668240031
transform 0 -1 2751 -1 0 -1058
box 0 0 2204 1138
use inv_buffer2  inv_buffer2_1
timestamp 1668240031
transform 0 1 5285 -1 0 -1058
box 0 0 2204 1138
use inv_buffer2  inv_buffer2_2
timestamp 1668240031
transform 0 -1 9326 -1 0 6219
box 0 0 2204 1138
use inv_buffer2  inv_buffer2_3
timestamp 1668240031
transform 0 1 -1289 -1 0 6230
box 0 0 2204 1138
use inv_simple1  inv_simple1_0
timestamp 1668240031
transform 0 -1 2138 1 0 6987
box -53 -613 858 525
use inv_simple1  inv_simple1_1
timestamp 1668240031
transform 0 1 3364 1 0 6987
box -53 -613 858 525
use inv_simple1  inv_simple1_2
timestamp 1668240031
transform 0 1 5898 1 0 6987
box -53 -613 858 525
use inv_simple1  inv_simple1_3
timestamp 1668240031
transform 0 -1 4672 1 0 6987
box -53 -613 858 525
use inv_simple1  inv_simple1_4
timestamp 1668240031
transform 0 -1 4672 -1 0 -201
box -53 -613 858 525
use inv_simple1  inv_simple1_5
timestamp 1668240031
transform 0 1 5898 -1 0 -201
box -53 -613 858 525
use inv_simple1  inv_simple1_6
timestamp 1668240031
transform 0 -1 2138 -1 0 -201
box -53 -613 858 525
use inv_simple1  inv_simple1_7
timestamp 1668240031
transform 0 1 3364 -1 0 -201
box -53 -613 858 525
use stf_ctrl  stf_ctrl_0
timestamp 1668240031
transform -1 0 12362 0 1 2267
box 1498 -2564 2762 3618
use vco_core_8  vco_core_8_0
timestamp 1668250571
transform 1 0 1484 0 1 4482
box -1484 -4482 6553 2304
<< labels >>
rlabel metal1 6511 -7137 6584 -7097 7 out2
port 1 n
rlabel metal1 4125 -7139 4198 -7099 7 out3
port 2 n
rlabel metal1 3842 -7139 3915 -7099 0 out4
port 3 n
rlabel metal1 1457 -7139 1530 -7099 3 out1
port 4 n
rlabel metal2 -1329 3363 -1200 3423 0 vdelay
port 5 n
rlabel metal1 8 2632 209 2832 0 vdd
port 6 n
rlabel metal1 379 2629 579 2829 6 vss
port 7 n
rlabel metal1 10780 771 10822 813 0 vbias
port 8 n
rlabel metal2 10822 1194 10864 1236 0 b0
port 9 n
rlabel metal2 10822 3240 10864 3282 0 b1
port 10 n
rlabel metal2 10822 5286 10864 5328 3 b2
port 11 n
rlabel metal1 3877 -4768 4163 -4671 7 vdd
rlabel metal1 3876 -5312 4162 -5215 3 vss
<< end >>
