magic
tech sky130A
magscale 1 2
timestamp 1668357910
<< pwell >>
rect -743 -280 743 280
<< nmos >>
rect -543 -70 -513 70
rect -447 -70 -417 70
rect -351 -70 -321 70
rect -255 -70 -225 70
rect -159 -70 -129 70
rect -63 -70 -33 70
rect 33 -70 63 70
rect 129 -70 159 70
rect 225 -70 255 70
rect 321 -70 351 70
rect 417 -70 447 70
rect 513 -70 543 70
<< ndiff >>
rect -609 58 -543 70
rect -609 -58 -593 58
rect -559 -58 -543 58
rect -609 -70 -543 -58
rect -513 58 -447 70
rect -513 -58 -497 58
rect -463 -58 -447 58
rect -513 -70 -447 -58
rect -417 58 -351 70
rect -417 -58 -401 58
rect -367 -58 -351 58
rect -417 -70 -351 -58
rect -321 58 -255 70
rect -321 -58 -305 58
rect -271 -58 -255 58
rect -321 -70 -255 -58
rect -225 58 -159 70
rect -225 -58 -209 58
rect -175 -58 -159 58
rect -225 -70 -159 -58
rect -129 58 -63 70
rect -129 -58 -113 58
rect -79 -58 -63 58
rect -129 -70 -63 -58
rect -33 58 33 70
rect -33 -58 -17 58
rect 17 -58 33 58
rect -33 -70 33 -58
rect 63 58 129 70
rect 63 -58 79 58
rect 113 -58 129 58
rect 63 -70 129 -58
rect 159 58 225 70
rect 159 -58 175 58
rect 209 -58 225 58
rect 159 -70 225 -58
rect 255 58 321 70
rect 255 -58 271 58
rect 305 -58 321 58
rect 255 -70 321 -58
rect 351 58 417 70
rect 351 -58 367 58
rect 401 -58 417 58
rect 351 -70 417 -58
rect 447 58 513 70
rect 447 -58 463 58
rect 497 -58 513 58
rect 447 -70 513 -58
rect 543 58 609 70
rect 543 -58 559 58
rect 593 -58 609 58
rect 543 -70 609 -58
<< ndiffc >>
rect -593 -58 -559 58
rect -497 -58 -463 58
rect -401 -58 -367 58
rect -305 -58 -271 58
rect -209 -58 -175 58
rect -113 -58 -79 58
rect -17 -58 17 58
rect 79 -58 113 58
rect 175 -58 209 58
rect 271 -58 305 58
rect 367 -58 401 58
rect 463 -58 497 58
rect 559 -58 593 58
<< psubdiff >>
rect -707 210 -611 244
rect 611 210 707 244
rect -707 148 -673 210
rect 673 148 707 210
rect -707 -210 -673 -148
rect 673 -210 707 -148
rect -707 -244 -611 -210
rect 611 -244 707 -210
<< psubdiffcont >>
rect -611 210 611 244
rect -707 -148 -673 148
rect 673 -148 707 148
rect -611 -244 611 -210
<< poly >>
rect -561 142 -495 158
rect -561 108 -545 142
rect -511 108 -495 142
rect -561 92 -495 108
rect 111 142 369 158
rect 111 108 127 142
rect 161 108 223 142
rect 257 108 319 142
rect 353 108 369 142
rect -543 70 -513 92
rect -447 70 -417 96
rect -351 70 -321 96
rect -255 70 -225 96
rect -159 70 -129 96
rect -63 70 -33 96
rect 33 70 63 96
rect 111 92 369 108
rect 495 142 561 158
rect 495 108 511 142
rect 545 108 561 142
rect 129 70 159 92
rect 225 70 255 92
rect 321 70 351 92
rect 417 70 447 96
rect 495 92 561 108
rect 513 70 543 92
rect -543 -96 -513 -70
rect -447 -92 -417 -70
rect -351 -92 -321 -70
rect -255 -92 -225 -70
rect -159 -92 -129 -70
rect -63 -92 -33 -70
rect 33 -92 63 -70
rect -465 -108 81 -92
rect 129 -96 159 -70
rect 225 -96 255 -70
rect 321 -96 351 -70
rect 417 -92 447 -70
rect -465 -142 -449 -108
rect -415 -142 -353 -108
rect -319 -142 -257 -108
rect -223 -142 -161 -108
rect -127 -142 -65 -108
rect -31 -142 31 -108
rect 65 -142 81 -108
rect -465 -158 81 -142
rect 399 -108 465 -92
rect 513 -96 543 -70
rect 399 -142 415 -108
rect 449 -142 465 -108
rect 399 -158 465 -142
<< polycont >>
rect -545 108 -511 142
rect 127 108 161 142
rect 223 108 257 142
rect 319 108 353 142
rect 511 108 545 142
rect -449 -142 -415 -108
rect -353 -142 -319 -108
rect -257 -142 -223 -108
rect -161 -142 -127 -108
rect -65 -142 -31 -108
rect 31 -142 65 -108
rect 415 -142 449 -108
<< locali >>
rect -707 210 -611 244
rect 611 210 707 244
rect -707 148 -673 210
rect -593 142 -559 210
rect 559 142 593 210
rect -593 108 -545 142
rect -511 108 -495 142
rect 111 108 127 142
rect 161 108 223 142
rect 257 108 319 142
rect 353 108 369 142
rect 495 108 511 142
rect 545 108 593 142
rect -593 58 -559 108
rect -593 -74 -559 -58
rect -497 58 -463 74
rect -497 -74 -463 -58
rect -401 58 -367 74
rect -401 -74 -367 -58
rect -305 58 -271 74
rect -305 -74 -271 -58
rect -209 58 -175 74
rect -209 -74 -175 -58
rect -113 58 -79 74
rect -113 -74 -79 -58
rect -17 58 17 74
rect -17 -74 17 -58
rect 79 58 113 74
rect 79 -74 113 -58
rect 175 58 209 74
rect 175 -74 209 -58
rect 271 58 305 74
rect 271 -74 305 -58
rect 367 58 401 74
rect 367 -74 401 -58
rect 463 58 497 74
rect 463 -74 497 -58
rect 559 58 593 108
rect 559 -74 593 -58
rect 673 148 707 210
rect -465 -142 -449 -108
rect -415 -142 -353 -108
rect -319 -142 -257 -108
rect -223 -142 -161 -108
rect -127 -142 -65 -108
rect -31 -142 31 -108
rect 65 -142 81 -108
rect 399 -142 415 -108
rect 449 -142 465 -108
rect -707 -210 -673 -148
rect 673 -210 707 -148
rect -707 -244 -611 -210
rect 611 -244 707 -210
<< viali >>
rect -545 108 -511 142
rect 127 108 161 142
rect 223 108 257 142
rect 319 108 353 142
rect 511 108 545 142
rect -593 -58 -559 58
rect -497 -58 -463 58
rect -401 -58 -367 58
rect -305 -58 -271 58
rect -209 -58 -175 58
rect -113 -58 -79 58
rect -17 -58 17 58
rect 79 -58 113 58
rect 175 -58 209 58
rect 271 -58 305 58
rect 367 -58 401 58
rect 463 -58 497 58
rect 559 -58 593 58
rect -449 -142 -415 -108
rect -353 -142 -319 -108
rect -257 -142 -223 -108
rect -161 -142 -127 -108
rect -65 -142 -31 -108
rect 31 -142 65 -108
rect 415 -142 449 -108
<< metal1 >>
rect -593 142 -499 148
rect -593 108 -545 142
rect -511 108 -499 142
rect -593 102 -499 108
rect 115 142 173 148
rect 211 142 269 148
rect 307 142 365 148
rect 115 108 127 142
rect 161 108 223 142
rect 257 108 319 142
rect 353 108 365 142
rect 115 102 173 108
rect 211 102 269 108
rect 307 102 365 108
rect 499 142 593 148
rect 499 108 511 142
rect 545 108 593 142
rect 499 102 593 108
rect -593 70 -557 102
rect 557 70 593 102
rect -599 58 -553 70
rect -599 0 -593 58
rect -609 -9 -593 0
rect -559 0 -553 58
rect -503 58 -457 70
rect -503 0 -497 58
rect -559 -9 -543 0
rect -609 -61 -602 -9
rect -550 -61 -543 -9
rect -609 -70 -543 -61
rect -513 -9 -497 0
rect -463 0 -457 58
rect -417 61 -351 70
rect -417 9 -410 61
rect -358 9 -351 61
rect -417 0 -401 9
rect -463 -9 -447 0
rect -513 -61 -506 -9
rect -454 -61 -447 -9
rect -513 -70 -447 -61
rect -407 -58 -401 0
rect -367 0 -351 9
rect -311 58 -265 70
rect -311 0 -305 58
rect -367 -58 -361 0
rect -407 -70 -361 -58
rect -321 -9 -305 0
rect -271 0 -265 58
rect -225 61 -159 70
rect -225 9 -218 61
rect -166 9 -159 61
rect -225 0 -209 9
rect -271 -9 -255 0
rect -321 -61 -314 -9
rect -262 -61 -255 -9
rect -321 -70 -255 -61
rect -215 -58 -209 0
rect -175 0 -159 9
rect -119 58 -73 70
rect -119 0 -113 58
rect -175 -58 -169 0
rect -215 -70 -169 -58
rect -129 -9 -113 0
rect -79 0 -73 58
rect -33 61 33 70
rect -33 9 -26 61
rect 26 9 33 61
rect -33 0 -17 9
rect -79 -9 -63 0
rect -129 -61 -122 -9
rect -70 -61 -63 -9
rect -129 -70 -63 -61
rect -23 -58 -17 0
rect 17 0 33 9
rect 73 58 119 70
rect 73 0 79 58
rect 17 -58 23 0
rect -23 -70 23 -58
rect 63 -9 79 0
rect 113 0 119 58
rect 159 61 225 70
rect 159 9 166 61
rect 218 9 225 61
rect 159 0 175 9
rect 113 -9 129 0
rect 63 -61 70 -9
rect 122 -61 129 -9
rect 63 -70 129 -61
rect 169 -58 175 0
rect 209 0 225 9
rect 265 58 311 70
rect 265 0 271 58
rect 209 -58 215 0
rect 169 -70 215 -58
rect 255 -9 271 0
rect 305 0 311 58
rect 351 61 417 70
rect 351 9 358 61
rect 410 9 417 61
rect 351 0 367 9
rect 305 -9 321 0
rect 255 -61 262 -9
rect 314 -61 321 -9
rect 255 -70 321 -61
rect 361 -58 367 0
rect 401 0 417 9
rect 457 58 503 70
rect 457 0 463 58
rect 401 -58 407 0
rect 361 -70 407 -58
rect 447 -9 463 0
rect 497 0 503 58
rect 553 58 599 70
rect 553 0 559 58
rect 497 -9 513 0
rect 447 -61 454 -9
rect 506 -61 513 -9
rect 447 -70 513 -61
rect 543 -9 559 0
rect 593 0 599 58
rect 593 -9 609 0
rect 543 -61 550 -9
rect 602 -61 609 -9
rect 543 -70 609 -61
rect -461 -108 -403 -102
rect -365 -108 -307 -102
rect -269 -108 -211 -102
rect -173 -108 -115 -102
rect -77 -108 -19 -102
rect 19 -108 77 -102
rect -461 -142 -449 -108
rect -415 -142 -353 -108
rect -319 -142 -257 -108
rect -223 -142 -161 -108
rect -127 -142 -65 -108
rect -31 -142 31 -108
rect 65 -142 77 -108
rect -461 -148 -403 -142
rect -365 -148 -307 -142
rect -269 -148 -211 -142
rect -173 -148 -115 -142
rect -77 -148 -19 -142
rect 19 -148 77 -142
rect 403 -108 461 -102
rect 403 -142 415 -108
rect 449 -142 495 -108
rect 403 -148 461 -142
<< via1 >>
rect -602 -58 -593 -9
rect -593 -58 -559 -9
rect -559 -58 -550 -9
rect -602 -61 -550 -58
rect -410 58 -358 61
rect -410 9 -401 58
rect -401 9 -367 58
rect -367 9 -358 58
rect -506 -58 -497 -9
rect -497 -58 -463 -9
rect -463 -58 -454 -9
rect -506 -61 -454 -58
rect -218 58 -166 61
rect -218 9 -209 58
rect -209 9 -175 58
rect -175 9 -166 58
rect -314 -58 -305 -9
rect -305 -58 -271 -9
rect -271 -58 -262 -9
rect -314 -61 -262 -58
rect -26 58 26 61
rect -26 9 -17 58
rect -17 9 17 58
rect 17 9 26 58
rect -122 -58 -113 -9
rect -113 -58 -79 -9
rect -79 -58 -70 -9
rect -122 -61 -70 -58
rect 166 58 218 61
rect 166 9 175 58
rect 175 9 209 58
rect 209 9 218 58
rect 70 -58 79 -9
rect 79 -58 113 -9
rect 113 -58 122 -9
rect 70 -61 122 -58
rect 358 58 410 61
rect 358 9 367 58
rect 367 9 401 58
rect 401 9 410 58
rect 262 -58 271 -9
rect 271 -58 305 -9
rect 305 -58 314 -9
rect 262 -61 314 -58
rect 454 -58 463 -9
rect 463 -58 497 -9
rect 497 -58 506 -9
rect 454 -61 506 -58
rect 550 -58 559 -9
rect 559 -58 593 -9
rect 593 -58 602 -9
rect 550 -61 602 -58
<< metal2 >>
rect -22 70 22 280
rect -417 61 417 70
rect -417 36 -410 61
rect -415 9 -410 36
rect -358 28 -218 61
rect -358 9 -353 28
rect -613 -8 -443 2
rect -415 0 -353 9
rect -223 9 -218 28
rect -166 28 -26 61
rect -166 9 -161 28
rect -223 0 -161 9
rect -31 9 -26 28
rect 26 28 166 61
rect 26 9 31 28
rect -31 0 31 9
rect 161 9 166 28
rect 218 28 358 61
rect 218 9 223 28
rect 161 0 223 9
rect 353 9 358 28
rect 410 36 417 61
rect 410 9 415 36
rect 353 0 415 9
rect -743 -9 -443 -8
rect -743 -50 -602 -9
rect -613 -61 -602 -50
rect -550 -61 -506 -9
rect -454 -28 -443 -9
rect -325 -9 -251 0
rect -325 -28 -314 -9
rect -454 -61 -314 -28
rect -262 -28 -251 -9
rect -133 -9 -59 0
rect -133 -28 -122 -9
rect -262 -61 -122 -28
rect -70 -28 -59 -9
rect 59 -9 133 0
rect 59 -28 70 -9
rect -70 -61 70 -28
rect 122 -28 133 -9
rect 251 -9 325 0
rect 251 -28 262 -9
rect 122 -61 262 -28
rect 314 -28 325 -9
rect 443 -8 613 2
rect 443 -9 743 -8
rect 443 -28 454 -9
rect 314 -61 454 -28
rect 506 -61 550 -9
rect 602 -50 743 -9
rect 602 -61 613 -50
rect -613 -70 613 -61
rect -613 -72 -443 -70
rect -325 -72 -251 -70
rect -133 -72 -59 -70
rect 59 -72 133 -70
rect 251 -72 325 -70
rect 443 -72 613 -70
<< labels >>
rlabel metal2 -22 234 22 278 7 in
port 1 n
rlabel metal2 -743 -50 -701 -8 1 vss
port 2 n
rlabel metal1 -17 -142 17 -108 0 swss
port 3 n
rlabel metal1 175 108 209 142 0 swtt
port 4 n
rlabel metal1 461 -142 495 -108 0 swff
port 5 n
<< properties >>
string FIXED_BBOX -690 -227 690 227
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.7 l 0.150 m 1 nf 12 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
