magic
tech sky130A
magscale 1 2
timestamp 1668153059
<< nwell >>
rect -455 -289 455 289
<< pmos >>
rect -255 -70 -225 70
rect -159 -70 -129 70
rect -63 -70 -33 70
rect 33 -70 63 70
rect 129 -70 159 70
rect 225 -70 255 70
<< pdiff >>
rect -317 58 -255 70
rect -317 -58 -305 58
rect -271 -58 -255 58
rect -317 -70 -255 -58
rect -225 58 -159 70
rect -225 -58 -209 58
rect -175 -58 -159 58
rect -225 -70 -159 -58
rect -129 58 -63 70
rect -129 -58 -113 58
rect -79 -58 -63 58
rect -129 -70 -63 -58
rect -33 58 33 70
rect -33 -58 -17 58
rect 17 -58 33 58
rect -33 -70 33 -58
rect 63 58 129 70
rect 63 -58 79 58
rect 113 -58 129 58
rect 63 -70 129 -58
rect 159 58 225 70
rect 159 -58 175 58
rect 209 -58 225 58
rect 159 -70 225 -58
rect 255 58 317 70
rect 255 -58 271 58
rect 305 -58 317 58
rect 255 -70 317 -58
<< pdiffc >>
rect -305 -58 -271 58
rect -209 -58 -175 58
rect -113 -58 -79 58
rect -17 -58 17 58
rect 79 -58 113 58
rect 175 -58 209 58
rect 271 -58 305 58
<< nsubdiff >>
rect -419 219 -323 253
rect 323 219 419 253
rect -419 157 -385 219
rect 385 157 419 219
rect -419 -219 -385 -157
rect 385 -219 419 -157
rect -419 -253 -323 -219
rect 323 -253 419 -219
<< nsubdiffcont >>
rect -323 219 323 253
rect -419 -157 -385 157
rect 385 -157 419 157
rect -323 -253 323 -219
<< poly >>
rect -273 151 -207 167
rect -273 117 -257 151
rect -223 117 -207 151
rect -273 101 -207 117
rect 207 151 273 167
rect 207 117 223 151
rect 257 117 273 151
rect 207 101 273 117
rect -255 70 -225 101
rect -159 70 -129 99
rect -63 70 -33 96
rect 33 70 63 99
rect 129 70 159 96
rect 225 70 255 101
rect -255 -96 -225 -70
rect -159 -101 -129 -70
rect -63 -101 -33 -70
rect 33 -101 63 -70
rect 129 -101 159 -70
rect 225 -96 255 -70
rect -177 -117 177 -101
rect -177 -151 -161 -117
rect -127 -151 -65 -117
rect -31 -151 31 -117
rect 65 -151 127 -117
rect 161 -151 177 -117
rect -177 -167 177 -151
<< polycont >>
rect -257 117 -223 151
rect 223 117 257 151
rect -161 -151 -127 -117
rect -65 -151 -31 -117
rect 31 -151 65 -117
rect 127 -151 161 -117
<< locali >>
rect -419 219 -323 253
rect 323 219 419 253
rect -419 157 -385 219
rect 385 157 419 219
rect -273 117 -257 151
rect -223 117 -207 151
rect 207 117 223 151
rect 257 117 273 151
rect -305 58 -271 74
rect -305 -74 -271 -58
rect -209 58 -175 74
rect -209 -74 -175 -58
rect -113 58 -79 74
rect -113 -74 -79 -58
rect -17 58 17 74
rect -17 -74 17 -58
rect 79 58 113 74
rect 79 -74 113 -58
rect 175 58 209 74
rect 175 -74 209 -58
rect 271 58 305 74
rect 271 -74 305 -58
rect -177 -151 -161 -117
rect -127 -151 -65 -117
rect -31 -151 31 -117
rect 65 -151 127 -117
rect 161 -151 177 -117
rect -419 -219 -385 -157
rect 385 -219 419 -157
rect -419 -253 -323 -219
rect 323 -253 419 -219
<< viali >>
rect -257 117 -223 151
rect 223 117 257 151
rect -305 -58 -271 58
rect -209 -58 -175 58
rect -113 -58 -79 58
rect -17 -58 17 58
rect 79 -58 113 58
rect 175 -58 209 58
rect 271 -58 305 58
rect -161 -151 -127 -117
rect -65 -151 -31 -117
rect 31 -151 65 -117
rect 127 -151 161 -117
<< metal1 >>
rect -305 151 -211 157
rect -305 117 -257 151
rect -223 117 -211 151
rect -305 111 -211 117
rect 211 151 305 157
rect 211 117 223 151
rect 257 117 305 151
rect 211 111 305 117
rect -305 70 -269 111
rect 269 70 305 111
rect -316 62 -164 70
rect -316 7 -314 62
rect -262 7 -218 62
rect -166 7 -164 62
rect -316 0 -305 7
rect -311 -58 -305 0
rect -271 0 -209 7
rect -271 -58 -265 0
rect -311 -70 -265 -58
rect -215 -58 -209 0
rect -175 0 -164 7
rect -119 58 -73 70
rect -119 0 -113 58
rect -175 -58 -169 0
rect -215 -70 -169 -58
rect -124 -7 -113 0
rect -79 0 -73 58
rect -28 62 28 70
rect -28 7 -26 62
rect 26 7 28 62
rect -28 0 -17 7
rect -79 -7 -68 0
rect -124 -62 -122 -7
rect -70 -62 -68 -7
rect -124 -70 -68 -62
rect -23 -58 -17 0
rect 17 0 28 7
rect 73 58 119 70
rect 73 0 79 58
rect 17 -58 23 0
rect -23 -70 23 -58
rect 68 -7 79 0
rect 113 0 119 58
rect 164 62 316 70
rect 164 7 166 62
rect 218 7 262 62
rect 314 7 316 62
rect 164 0 175 7
rect 113 -7 124 0
rect 68 -62 70 -7
rect 122 -62 124 -7
rect 68 -70 124 -62
rect 169 -58 175 0
rect 209 0 271 7
rect 209 -58 215 0
rect 169 -70 215 -58
rect 265 -58 271 0
rect 305 0 316 7
rect 305 -58 311 0
rect 265 -70 311 -58
rect -173 -117 -115 -111
rect -77 -117 -19 -111
rect 19 -117 77 -111
rect 115 -117 173 -111
rect -177 -151 -161 -117
rect -127 -151 -65 -117
rect -31 -151 31 -117
rect 65 -151 127 -117
rect 161 -151 177 -117
rect -173 -157 -115 -151
rect -77 -157 -19 -151
rect 19 -157 77 -151
rect 115 -157 173 -151
<< via1 >>
rect -314 58 -262 62
rect -314 7 -305 58
rect -305 7 -271 58
rect -271 7 -262 58
rect -218 58 -166 62
rect -218 7 -209 58
rect -209 7 -175 58
rect -175 7 -166 58
rect -26 58 26 62
rect -26 7 -17 58
rect -17 7 17 58
rect 17 7 26 58
rect -122 -58 -113 -7
rect -113 -58 -79 -7
rect -79 -58 -70 -7
rect -122 -62 -70 -58
rect 166 58 218 62
rect 166 7 175 58
rect 175 7 209 58
rect 209 7 218 58
rect 262 58 314 62
rect 262 7 271 58
rect 271 7 305 58
rect 305 7 314 58
rect 70 -58 79 -7
rect 79 -58 113 -7
rect 113 -58 122 -7
rect 70 -62 122 -58
<< metal2 >>
rect -316 62 316 70
rect -316 7 -314 62
rect -262 7 -218 62
rect -166 28 -26 62
rect -166 7 -164 28
rect -316 0 -164 7
rect -28 7 -26 28
rect 26 28 166 62
rect 26 7 28 28
rect -28 0 28 7
rect 164 7 166 28
rect 218 7 262 62
rect 314 7 316 62
rect 164 0 316 7
rect -124 -7 -68 0
rect -124 -62 -122 -7
rect -70 -28 -68 -7
rect 68 -7 124 0
rect 68 -28 70 -7
rect -70 -62 70 -28
rect 122 -62 124 -7
rect -124 -70 124 -62
<< properties >>
string FIXED_BBOX -402 -236 402 236
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.7 l 0.15 m 1 nf 6 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
