magic
tech sky130A
magscale 1 2
timestamp 1668163051
<< metal2 >>
rect 73442 12503 74458 12600
rect 73440 12331 74458 12503
rect 71224 10791 71794 11361
rect 73440 11215 73658 12331
rect 74253 11215 74458 12331
rect 73440 10942 74458 11215
<< via2 >>
rect 73658 11215 74253 12331
<< metal3 >>
rect 73440 12331 74458 19661
rect 73440 11215 73658 12331
rect 74253 11215 74458 12331
rect 73440 10942 74458 11215
use cap_200p  cap_200p_0
timestamp 1668108937
transform 1 0 44238 0 1 22632
box -3186 -3040 60524 67041
use r_8k  r_8k_1
timestamp 1668153059
transform 1 0 72736 0 1 8422
box -2496 -2369 2460 2830
<< end >>
