magic
tech sky130A
magscale 1 2
timestamp 1659939748
<< error_p >>
rect -269 -108 -211 -102
rect 211 -108 269 -102
rect -269 -142 -257 -108
rect 211 -142 223 -108
rect -269 -148 -211 -142
rect 211 -148 269 -142
<< pwell >>
rect -455 -280 455 280
<< nmos >>
rect -255 -70 -225 70
rect -159 -70 -129 70
rect -63 -70 -33 70
rect 33 -70 63 70
rect 129 -70 159 70
rect 225 -70 255 70
<< ndiff >>
rect -325 58 -255 70
rect -325 -2 -305 58
rect -317 -58 -305 -2
rect -271 -58 -255 58
rect -317 -70 -255 -58
rect -225 58 -159 70
rect -225 -58 -209 58
rect -175 -58 -159 58
rect -225 -70 -159 -58
rect -129 58 -63 70
rect -129 -58 -113 58
rect -79 -58 -63 58
rect -129 -70 -63 -58
rect -33 58 33 70
rect -33 -58 -17 58
rect 17 -58 33 58
rect -33 -70 33 -58
rect 63 58 129 70
rect 63 -58 79 58
rect 113 -58 129 58
rect 63 -70 129 -58
rect 159 58 225 70
rect 159 -58 175 58
rect 209 -58 225 58
rect 159 -70 225 -58
rect 255 58 325 70
rect 255 -58 271 58
rect 305 -2 325 58
rect 305 -58 317 -2
rect 255 -70 317 -58
<< ndiffc >>
rect -305 -58 -271 58
rect -209 -58 -175 58
rect -113 -58 -79 58
rect -17 -58 17 58
rect 79 -58 113 58
rect 175 -58 209 58
rect 271 -58 305 58
<< psubdiff >>
rect -419 210 -323 244
rect 323 210 419 244
rect -419 148 -385 210
rect 385 148 419 210
rect -419 -210 -385 -148
rect 385 -210 419 -148
rect -419 -244 -323 -210
rect 323 -244 419 -210
<< psubdiffcont >>
rect -323 210 323 244
rect -419 -148 -385 148
rect 385 -148 419 148
rect -323 -244 323 -210
<< poly >>
rect -177 142 177 158
rect -177 108 -161 142
rect -127 108 -65 142
rect -31 108 31 142
rect 65 108 127 142
rect 161 108 177 142
rect -255 70 -225 96
rect -177 92 177 108
rect -159 70 -129 92
rect -63 70 -33 92
rect 33 70 63 92
rect 129 70 159 92
rect 225 70 255 96
rect -255 -92 -225 -70
rect -273 -108 -207 -92
rect -159 -96 -129 -70
rect -63 -96 -33 -70
rect 33 -96 63 -70
rect 129 -96 159 -70
rect 225 -92 255 -70
rect -273 -142 -257 -108
rect -223 -142 -207 -108
rect -273 -158 -207 -142
rect 207 -108 273 -92
rect 207 -142 223 -108
rect 257 -142 273 -108
rect 207 -158 273 -142
<< polycont >>
rect -161 108 -127 142
rect -65 108 -31 142
rect 31 108 65 142
rect 127 108 161 142
rect -257 -142 -223 -108
rect 223 -142 257 -108
<< locali >>
rect -419 210 -323 244
rect 323 210 419 244
rect -419 148 -385 210
rect -525 -1 -455 69
rect 385 148 419 210
rect -177 108 -161 142
rect -127 108 -65 142
rect -31 108 31 142
rect 65 108 127 142
rect 161 108 177 142
rect -305 58 -271 74
rect -305 -74 -271 -58
rect -209 58 -175 74
rect -209 -74 -175 -58
rect -113 58 -79 74
rect -113 -74 -79 -58
rect -17 58 17 74
rect -17 -74 17 -58
rect 79 58 113 74
rect 79 -74 113 -58
rect 175 58 209 74
rect 175 -74 209 -58
rect 271 58 305 74
rect 271 -74 305 -58
rect -273 -142 -257 -108
rect -223 -142 -207 -108
rect 207 -142 223 -108
rect 257 -142 273 -108
rect -419 -210 -385 -148
rect 385 -210 419 -148
rect -419 -244 -323 -210
rect 323 -244 419 -210
<< viali >>
rect -161 108 -127 142
rect -65 108 -31 142
rect 31 108 65 142
rect 127 108 161 142
rect -305 -58 -271 58
rect -209 -58 -175 58
rect -113 -58 -79 58
rect -17 -58 17 58
rect 79 -58 113 58
rect 175 -58 209 58
rect 271 -58 305 58
rect -257 -142 -223 -108
rect 223 -142 257 -108
<< metal1 >>
rect -173 142 -115 148
rect -77 142 -19 148
rect 19 142 77 148
rect 115 142 173 148
rect -173 108 -161 142
rect -127 108 -65 142
rect -31 108 31 142
rect 65 108 127 142
rect 161 108 173 142
rect -173 102 -115 108
rect -77 102 -19 108
rect 19 102 77 108
rect 115 102 173 108
rect -318 61 -258 70
rect -318 9 -314 61
rect -262 9 -258 61
rect -318 0 -305 9
rect -311 -58 -305 0
rect -271 0 -258 9
rect -222 61 -162 70
rect -222 9 -218 61
rect -166 9 -162 61
rect -222 0 -209 9
rect -271 -58 -265 0
rect -311 -70 -265 -58
rect -215 -58 -209 0
rect -175 0 -162 9
rect -119 58 -73 70
rect -119 0 -113 58
rect -175 -58 -169 0
rect -215 -70 -169 -58
rect -126 -9 -113 0
rect -79 0 -73 58
rect -30 61 30 70
rect -30 9 -26 61
rect 26 9 30 61
rect -30 0 -17 9
rect -79 -9 -66 0
rect -126 -61 -122 -9
rect -70 -61 -66 -9
rect -126 -70 -66 -61
rect -23 -58 -17 0
rect 17 0 30 9
rect 73 58 119 70
rect 73 0 79 58
rect 17 -58 23 0
rect -23 -70 23 -58
rect 66 -9 79 0
rect 113 0 119 58
rect 162 61 222 70
rect 162 9 166 61
rect 218 9 222 61
rect 162 0 175 9
rect 113 -9 126 0
rect 66 -61 70 -9
rect 122 -61 126 -9
rect 66 -70 126 -61
rect 169 -58 175 0
rect 209 0 222 9
rect 258 61 318 70
rect 258 9 262 61
rect 314 9 318 61
rect 258 0 271 9
rect 209 -58 215 0
rect 169 -70 215 -58
rect 265 -58 271 0
rect 305 0 318 9
rect 305 -58 311 0
rect 265 -70 311 -58
rect -269 -108 -211 -102
rect -269 -142 -257 -108
rect -223 -142 -211 -108
rect -269 -148 -211 -142
rect 211 -108 269 -102
rect 211 -142 223 -108
rect 257 -142 269 -108
rect 211 -148 269 -142
<< via1 >>
rect -314 58 -262 61
rect -314 9 -305 58
rect -305 9 -271 58
rect -271 9 -262 58
rect -218 58 -166 61
rect -218 9 -209 58
rect -209 9 -175 58
rect -175 9 -166 58
rect -26 58 26 61
rect -26 9 -17 58
rect -17 9 17 58
rect 17 9 26 58
rect -122 -58 -113 -9
rect -113 -58 -79 -9
rect -79 -58 -70 -9
rect -122 -61 -70 -58
rect 166 58 218 61
rect 166 9 175 58
rect 175 9 209 58
rect 209 9 218 58
rect 70 -58 79 -9
rect 79 -58 113 -9
rect 113 -58 122 -9
rect 70 -61 122 -58
rect 262 58 314 61
rect 262 9 271 58
rect 271 9 305 58
rect 305 9 314 58
<< metal2 >>
rect -325 63 -155 72
rect -325 7 -316 63
rect -260 7 -220 63
rect -164 7 -155 63
rect -325 -2 -155 7
rect -37 63 37 72
rect -37 7 -28 63
rect 28 7 37 63
rect -126 -9 -66 0
rect -37 -2 37 7
rect 155 63 325 72
rect 155 7 164 63
rect 220 7 260 63
rect 316 7 325 63
rect -126 -61 -122 -9
rect -70 -36 -66 -9
rect 66 -9 126 0
rect 155 -2 325 7
rect 66 -36 70 -9
rect -70 -61 70 -36
rect 122 -36 126 -9
rect 122 -61 129 -36
rect -126 -70 129 -61
<< via2 >>
rect -316 61 -260 63
rect -316 9 -314 61
rect -314 9 -262 61
rect -262 9 -260 61
rect -316 7 -260 9
rect -220 61 -164 63
rect -220 9 -218 61
rect -218 9 -166 61
rect -166 9 -164 61
rect -220 7 -164 9
rect -28 61 28 63
rect -28 9 -26 61
rect -26 9 26 61
rect 26 9 28 61
rect -28 7 28 9
rect 164 61 220 63
rect 164 9 166 61
rect 166 9 218 61
rect 218 9 220 61
rect 164 7 220 9
rect 260 61 316 63
rect 260 9 262 61
rect 262 9 314 61
rect 314 9 316 61
rect 260 7 316 9
<< metal3 >>
rect -325 70 -155 72
rect -37 70 37 72
rect 155 70 325 72
rect -325 63 325 70
rect -325 7 -316 63
rect -260 7 -220 63
rect -164 10 -28 63
rect -164 7 -155 10
rect -325 -2 -155 7
rect -37 7 -28 10
rect 28 10 164 63
rect 28 7 37 10
rect -37 -2 37 7
rect 155 7 164 10
rect 220 7 260 63
rect 316 7 325 63
rect 155 -2 325 7
<< properties >>
string FIXED_BBOX -402 -227 402 227
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.7 l 0.150 m 1 nf 6 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
