magic
tech sky130A
magscale 1 2
timestamp 1668153059
<< metal1 >>
rect 514 958 578 964
rect 514 950 520 958
rect 508 916 520 950
rect 514 906 520 916
rect 572 906 578 958
rect 514 900 578 906
rect 226 686 290 692
rect 226 634 232 686
rect 284 678 290 686
rect 284 644 296 678
rect 284 634 290 644
rect 226 628 290 634
rect 226 532 290 538
rect 226 480 232 532
rect 284 524 290 532
rect 514 532 578 538
rect 514 524 520 532
rect 284 490 323 524
rect 481 490 520 524
rect 284 480 289 490
rect 226 471 289 480
rect 514 480 520 490
rect 572 480 578 532
rect 514 474 578 480
rect -537 437 289 471
rect 515 471 578 474
rect 515 437 1341 471
rect -1147 297 -1111 375
rect -245 -53 -211 437
rect -175 403 -123 409
rect -175 345 -123 351
rect 927 403 979 409
rect 927 345 979 351
rect -315 -87 -211 -53
rect -315 -99 -266 -87
rect -166 -99 -132 345
rect -87 85 232 119
rect 572 85 891 119
rect -87 -53 -53 85
rect 857 -53 891 85
rect -87 -87 16 -53
rect -33 -99 16 -87
rect 787 -87 891 -53
rect 787 -99 836 -87
rect 936 -99 970 345
rect 1015 -53 1049 437
rect 1015 -87 1118 -53
rect 1069 -99 1118 -87
rect -330 -105 -266 -99
rect -330 -157 -324 -105
rect -272 -157 -266 -105
rect -330 -163 -266 -157
rect -182 -105 -118 -99
rect -182 -157 -176 -105
rect -124 -157 -118 -105
rect -182 -163 -118 -157
rect -33 -105 31 -99
rect -33 -157 -27 -105
rect 25 -157 31 -105
rect -33 -163 31 -157
rect 772 -105 836 -99
rect 772 -157 778 -105
rect 830 -157 836 -105
rect 772 -163 836 -157
rect 920 -105 984 -99
rect 920 -157 926 -105
rect 978 -157 984 -105
rect 920 -163 984 -157
rect 1069 -105 1133 -99
rect 1069 -157 1075 -105
rect 1127 -157 1133 -105
rect 1069 -163 1133 -157
rect -730 -234 -724 -182
rect -672 -234 -666 -182
rect 1470 -234 1476 -182
rect 1528 -234 1534 -182
rect -719 -364 -677 -234
rect 610 -325 616 -273
rect 668 -325 674 -273
rect 1481 -364 1523 -234
rect -730 -416 -724 -364
rect -672 -416 -666 -364
rect 1470 -416 1476 -364
rect 1528 -416 1534 -364
rect 1145 -563 1151 -554
rect 863 -597 1151 -563
rect 433 -665 467 -597
rect 1145 -606 1151 -597
rect 1203 -606 1209 -554
rect 1145 -665 1151 -656
rect 433 -699 1151 -665
rect 1145 -708 1151 -699
rect 1203 -708 1209 -656
<< via1 >>
rect 520 906 572 958
rect 232 634 284 686
rect 232 480 284 532
rect 520 480 572 532
rect -175 351 -123 403
rect 927 351 979 403
rect -324 -157 -272 -105
rect -176 -157 -124 -105
rect -27 -157 25 -105
rect 778 -157 830 -105
rect 926 -157 978 -105
rect 1075 -157 1127 -105
rect -724 -234 -672 -182
rect 1476 -234 1528 -182
rect 616 -325 668 -273
rect -724 -416 -672 -364
rect 1476 -416 1528 -364
rect 1151 -606 1203 -554
rect 1151 -708 1203 -656
<< metal2 >>
rect 385 1049 419 1085
rect -115 1015 919 1049
rect 508 960 584 970
rect 508 904 518 960
rect 574 904 584 960
rect 508 894 584 904
rect 220 688 296 698
rect 220 632 230 688
rect 286 632 296 688
rect 220 622 296 632
rect 220 534 296 544
rect 220 478 230 534
rect 286 478 296 534
rect -489 437 -132 471
rect 220 468 296 478
rect 508 534 584 544
rect 508 478 518 534
rect 574 478 584 534
rect 508 468 584 478
rect -166 403 -132 437
rect 936 437 1293 471
rect 936 403 970 437
rect -181 351 -175 403
rect -123 351 -117 403
rect 921 351 927 403
rect 979 351 985 403
rect 936 349 970 351
rect -719 -176 -677 157
rect -335 -103 -261 -94
rect -335 -159 -326 -103
rect -270 -159 -261 -103
rect -335 -168 -261 -159
rect -188 -103 -112 -93
rect -188 -159 -178 -103
rect -122 -159 -112 -103
rect -188 -169 -112 -159
rect -38 -103 36 -94
rect -38 -159 -29 -103
rect 27 -159 36 -103
rect -38 -168 36 -159
rect 380 -175 424 157
rect 767 -103 841 -94
rect 767 -159 776 -103
rect 832 -159 841 -103
rect 767 -168 841 -159
rect 914 -103 990 -93
rect 914 -159 924 -103
rect 980 -159 990 -103
rect 914 -169 990 -159
rect 1064 -103 1138 -94
rect 1064 -159 1073 -103
rect 1129 -159 1138 -103
rect 1064 -168 1138 -159
rect 1481 -176 1523 157
rect -724 -182 -672 -176
rect -724 -240 -672 -234
rect 1476 -182 1528 -176
rect 1476 -240 1528 -234
rect 616 -273 668 -267
rect 668 -316 1669 -282
rect 616 -331 668 -325
rect -724 -364 -672 -358
rect -724 -422 -672 -416
rect 1476 -364 1528 -358
rect 1476 -422 1528 -416
rect -719 -463 -677 -422
rect 1481 -463 1523 -422
rect -719 -505 -341 -463
rect 1145 -505 1523 -463
rect 1151 -554 1203 -548
rect 1203 -597 1669 -563
rect 1151 -612 1203 -606
rect 1151 -656 1203 -650
rect 1203 -699 1669 -665
rect 1151 -714 1203 -708
<< via2 >>
rect 518 958 574 960
rect 518 906 520 958
rect 520 906 572 958
rect 572 906 574 958
rect 518 904 574 906
rect 230 686 286 688
rect 230 634 232 686
rect 232 634 284 686
rect 284 634 286 686
rect 230 632 286 634
rect 230 532 286 534
rect 230 480 232 532
rect 232 480 284 532
rect 284 480 286 532
rect 230 478 286 480
rect 518 532 574 534
rect 518 480 520 532
rect 520 480 572 532
rect 572 480 574 532
rect 518 478 574 480
rect -326 -105 -270 -103
rect -326 -157 -324 -105
rect -324 -157 -272 -105
rect -272 -157 -270 -105
rect -326 -159 -270 -157
rect -178 -105 -122 -103
rect -178 -157 -176 -105
rect -176 -157 -124 -105
rect -124 -157 -122 -105
rect -178 -159 -122 -157
rect -29 -105 27 -103
rect -29 -157 -27 -105
rect -27 -157 25 -105
rect 25 -157 27 -105
rect -29 -159 27 -157
rect 776 -105 832 -103
rect 776 -157 778 -105
rect 778 -157 830 -105
rect 830 -157 832 -105
rect 776 -159 832 -157
rect 924 -105 980 -103
rect 924 -157 926 -105
rect 926 -157 978 -105
rect 978 -157 980 -105
rect 924 -159 980 -157
rect 1073 -105 1129 -103
rect 1073 -157 1075 -105
rect 1075 -157 1127 -105
rect 1127 -157 1129 -105
rect 1073 -159 1129 -157
<< metal3 >>
rect 502 964 590 976
rect 502 900 514 964
rect 578 962 590 964
rect 578 902 621 962
rect 578 900 590 902
rect 502 888 590 900
rect -1581 805 -1450 865
rect -998 805 -732 865
rect -280 805 -11 865
rect 815 805 1084 865
rect 1536 805 1669 865
rect 214 692 302 704
rect 214 690 226 692
rect 183 630 226 690
rect 214 628 226 630
rect 290 628 302 692
rect 214 616 302 628
rect 214 538 302 550
rect 214 536 226 538
rect 183 476 226 536
rect 214 474 226 476
rect 290 474 302 538
rect 214 462 302 474
rect 502 538 590 550
rect 502 474 514 538
rect 578 536 590 538
rect 578 476 621 536
rect 578 474 590 476
rect 502 462 590 474
rect -1581 157 -1354 217
rect -998 157 -732 217
rect -376 157 1180 217
rect 1536 157 1669 217
rect -179 -87 -119 -56
rect 923 -87 983 -56
rect -335 -103 -261 -94
rect -335 -159 -326 -103
rect -270 -159 -261 -103
rect -335 -168 -261 -159
rect -194 -99 -106 -87
rect -194 -163 -182 -99
rect -118 -163 -106 -99
rect -328 -245 -268 -168
rect -194 -175 -106 -163
rect -38 -103 36 -94
rect -38 -159 -29 -103
rect 27 -159 36 -103
rect -38 -168 36 -159
rect 767 -103 841 -94
rect 767 -159 776 -103
rect 832 -159 841 -103
rect 767 -168 841 -159
rect 908 -99 996 -87
rect 908 -163 920 -99
rect 984 -163 996 -99
rect -31 -245 29 -168
rect 774 -245 834 -168
rect 908 -175 996 -163
rect 1064 -103 1138 -94
rect 1064 -159 1073 -103
rect 1129 -159 1138 -103
rect 1064 -168 1138 -159
rect 1071 -245 1131 -168
<< via3 >>
rect 514 960 578 964
rect 514 904 518 960
rect 518 904 574 960
rect 574 904 578 960
rect 514 900 578 904
rect 226 688 290 692
rect 226 632 230 688
rect 230 632 286 688
rect 286 632 290 688
rect 226 628 290 632
rect 226 534 290 538
rect 226 478 230 534
rect 230 478 286 534
rect 286 478 290 534
rect 226 474 290 478
rect 514 534 578 538
rect 514 478 518 534
rect 518 478 574 534
rect 574 478 578 534
rect 514 474 578 478
rect -182 -103 -118 -99
rect -182 -159 -178 -103
rect -178 -159 -122 -103
rect -122 -159 -118 -103
rect -182 -163 -118 -159
rect 920 -103 984 -99
rect 920 -159 924 -103
rect 924 -159 980 -103
rect 980 -159 984 -103
rect 920 -163 984 -159
<< metal4 >>
rect -179 -87 -119 1083
rect 228 704 288 1083
rect 516 976 576 1083
rect 502 964 590 976
rect 502 900 514 964
rect 578 900 590 964
rect 502 888 590 900
rect 214 692 302 704
rect 214 628 226 692
rect 290 628 302 692
rect 214 616 302 628
rect 228 550 288 616
rect 516 550 576 888
rect 214 538 302 550
rect 214 474 226 538
rect 290 474 302 538
rect 214 462 302 474
rect 502 538 590 550
rect 502 474 514 538
rect 578 474 590 538
rect 502 462 590 474
rect 923 -87 983 1083
rect -194 -99 -106 -87
rect -194 -163 -182 -99
rect -118 -163 -106 -99
rect -194 -175 -106 -163
rect 908 -99 996 -87
rect 908 -163 920 -99
rect 984 -163 996 -99
rect 908 -175 996 -163
use current_tails_1  current_tails_1_0
timestamp 1668153059
transform 1 0 402 0 1 -455
box -743 -280 743 280
use n_cell_3  n_cell_3_0
timestamp 1668153059
transform -1 0 -1175 0 1 227
box -310 -280 310 280
use n_cell_3  sky130_fd_pr__nfet_01v8_5ZA63U_0
timestamp 1668153059
transform 1 0 -555 0 1 227
box -310 -280 310 280
use n_cell_3  sky130_fd_pr__nfet_01v8_5ZA63U_1
timestamp 1668153059
transform -1 0 1359 0 1 227
box -310 -280 310 280
use n_cell_1  sky130_fd_pr__nfet_01v8_lvt_GVQ53W_0
timestamp 1668153059
transform 1 0 402 0 1 227
box -455 -280 455 280
use p_cell_3  sky130_fd_pr__pfet_01v8_X6PFBL_0
timestamp 1668153059
transform 1 0 402 0 1 796
box -551 -289 551 289
use sky130_fd_pr__pfet_01v8_X679XQ  sky130_fd_pr__pfet_01v8_X679XQ_0
timestamp 1668153059
transform 1 0 -507 0 -1 795
box -358 -288 358 288
use sky130_fd_pr__pfet_01v8_X679XQ  sky130_fd_pr__pfet_01v8_X679XQ_1
timestamp 1668153059
transform -1 0 1311 0 -1 795
box -358 -288 358 288
use sky130_fd_pr__pfet_01v8_X679XQ  sky130_fd_pr__pfet_01v8_X679XQ_2
timestamp 1668153059
transform -1 0 -1223 0 -1 795
box -358 -288 358 288
<< labels >>
rlabel metal1 -87 -87 -53 -53 0 din1
port 1 n
rlabel metal1 857 -87 891 -53 5 din2
port 2 n
rlabel metal3 -1581 805 -1521 865 0 vdd
port 4 n
rlabel metal1 -53 437 -19 471 4 dout1
port 5 n
rlabel metal1 823 437 857 471 3 dout2
port 6 n
rlabel metal2 385 1015 419 1085 4 vb
port 7 n
rlabel metal2 1635 -316 1669 -282 3 b1
port 8 n
rlabel metal2 1635 -597 1669 -563 6 b0
port 9 n
rlabel metal2 1635 -699 1669 -665 0 b2
port 10 n
rlabel metal2 380 -122 424 -78 3 net1
rlabel metal3 -1581 157 -1521 217 0 vss
port 3 n
<< end >>
