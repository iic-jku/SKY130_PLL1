magic
tech sky130A
magscale 1 2
timestamp 1661285251
<< metal1 >>
rect 3808 3710 3814 3762
rect 3866 3710 3872 3762
rect 3687 3679 3721 3685
rect 3672 3627 3678 3679
rect 3730 3627 3736 3679
rect 3687 3621 3721 3627
rect 3551 3596 3585 3602
rect 3536 3544 3542 3596
rect 3594 3544 3600 3596
rect 3551 3538 3585 3544
<< via1 >>
rect 3814 3710 3866 3762
rect 3678 3627 3730 3679
rect 3542 3544 3594 3596
<< metal2 >>
rect 2420 5787 2454 6846
rect 4954 5764 4988 6918
rect 10297 5779 10339 5821
rect 12345 5779 12387 5821
rect 14393 5779 14435 5821
rect 7482 5425 7491 5485
rect 7551 5476 7560 5485
rect 7551 5434 7704 5476
rect 7551 5425 7560 5434
rect 7482 4777 7491 4837
rect 7551 4828 7560 4837
rect 7551 4809 7844 4828
rect 7551 4786 7896 4809
rect 7551 4777 7560 4786
rect 7802 4767 7896 4786
rect 3814 3762 3866 3768
rect 10297 3753 10339 4515
rect 3866 3719 10339 3753
rect 3814 3704 3866 3710
rect 3678 3679 3730 3685
rect 12345 3670 12387 4515
rect 3730 3636 12387 3670
rect 3678 3621 3730 3627
rect 3542 3596 3594 3602
rect 14393 3587 14435 4515
rect 3594 3553 14435 3587
rect 3542 3538 3594 3544
<< via2 >>
rect 7491 5425 7551 5485
rect 7491 4777 7551 4837
<< metal3 >>
rect 7486 5485 7556 5490
rect 6298 5425 7491 5485
rect 7551 5425 7556 5485
rect 7486 5420 7556 5425
rect 7486 4837 7556 4842
rect 6298 4777 7491 4837
rect 7551 4777 7556 4837
rect 7486 4772 7556 4777
<< metal4 >>
rect 1856 5763 1916 6846
rect 2958 5760 3018 6846
rect 6238 4273 7468 4333
rect 6238 4013 7468 4073
rect 6238 3753 6298 3813
rect 6238 3493 6298 3553
rect 6238 3233 6298 3293
rect 6238 2973 6298 3033
rect 6238 2713 6298 2773
rect 6238 2453 6298 2513
use stf_ctrl  stf_ctrl_0 ma2022
timestamp 1661273666
transform 0 1 11374 -1 0 7277
box 1498 -3670 2762 3618
use vco_core_8  vco_core_8_0 ma2022
timestamp 1661242302
transform 1 0 1170 0 1 4482
box -1170 -4482 6238 2304
<< labels >>
rlabel metal2 7408 3719 7442 3753 5 b0
rlabel metal2 7408 3636 7442 3670 0 b1
rlabel metal2 7408 3553 7442 3587 5 b2
rlabel metal3 7408 4777 7468 4837 3 vss
rlabel metal3 7408 5425 7468 5485 3 vdd
rlabel metal2 2420 6786 2454 6820 4 vb2
rlabel metal2 4954 6786 4988 6820 0 vb1
rlabel metal4 7408 4013 7468 4073 0 out2
rlabel metal4 7408 4273 7468 4333 0 out1
rlabel metal4 1856 6786 1916 6846 8 inv1
rlabel metal4 2958 6786 3018 6846 0 inv2
<< end >>
