magic
tech sky130A
magscale 1 2
timestamp 1669727735
<< metal1 >>
rect -2272 3139 -1422 3145
rect -2272 1622 -1422 2289
rect 2138 3139 2988 3145
rect 2138 1622 2988 2289
rect -2252 -938 -1432 -138
rect 2158 -936 2978 -136
rect -2232 -1770 -1432 -938
rect -2232 -2576 -1432 -2570
rect 2178 -1768 2978 -936
rect 2178 -2574 2978 -2568
<< via1 >>
rect -2272 2289 -1422 3139
rect 2138 2289 2988 3139
rect -2245 41 -1451 644
rect 2163 38 2960 647
rect -2232 -2570 -1432 -1770
rect 2178 -2568 2978 -1768
<< metal2 >>
rect -2272 3139 -1422 3148
rect -2278 2289 -2272 3139
rect -1422 2289 -1416 3139
rect -999 2731 567 3372
rect 2138 3139 2988 3148
rect -2272 2280 -1422 2289
rect -999 662 -359 2731
rect 2132 2289 2138 3139
rect 2988 2289 2994 3139
rect 2138 2280 2988 2289
rect -2262 644 -359 662
rect -2262 41 -2245 644
rect -1451 41 -359 644
rect 168 647 2978 662
rect 168 89 2163 647
rect -2262 22 -359 41
rect 169 38 2163 89
rect 2960 38 2978 647
rect 169 22 2978 38
rect -2252 -938 -1432 -138
rect 2158 -936 2978 -136
rect -2232 -1770 -1432 -1761
rect 2178 -1768 2978 -1759
rect -2238 -2570 -2232 -1770
rect -1432 -2570 -1426 -1770
rect 2172 -2568 2178 -1768
rect 2978 -2568 2984 -1768
rect -2232 -2579 -1432 -2570
rect 2178 -2577 2978 -2568
<< via2 >>
rect -2272 2289 -1422 3139
rect 2138 2289 2988 3139
rect -2232 -2570 -1432 -1770
rect 2178 -2568 2978 -1768
<< metal3 >>
rect -2277 3144 -1417 3150
rect -2277 2289 -2272 2294
rect -1422 2289 -1417 2294
rect -2277 2284 -1417 2289
rect 2133 3144 2993 3150
rect 2133 2289 2138 2294
rect 2988 2289 2993 2294
rect 2133 2284 2993 2289
rect -2237 -1770 -1427 -1765
rect -2237 -1775 -2232 -1770
rect -1432 -1775 -1427 -1770
rect -2237 -2581 -1427 -2575
rect 2173 -1768 2983 -1763
rect 2173 -1773 2178 -1768
rect 2978 -1773 2983 -1768
rect 2173 -2579 2983 -2573
<< via3 >>
rect -2277 3139 -1417 3144
rect -2277 2294 -2272 3139
rect -2272 2294 -1422 3139
rect -1422 2294 -1417 3139
rect 2133 3139 2993 3144
rect 2133 2294 2138 3139
rect 2138 2294 2988 3139
rect 2988 2294 2993 3139
rect -2237 -2570 -2232 -1775
rect -2232 -2570 -1432 -1775
rect -1432 -2570 -1427 -1775
rect -2237 -2575 -1427 -2570
rect 2173 -2568 2178 -1773
rect 2178 -2568 2978 -1773
rect 2978 -2568 2983 -1773
rect 2173 -2573 2983 -2568
<< metal4 >>
rect -2278 2294 -2277 2295
rect -1417 2294 -1416 2295
rect -2278 2293 -1416 2294
rect 2132 2294 2133 2295
rect 2993 2294 2994 2295
rect 2132 2293 2994 2294
rect 2172 -1773 2984 -1772
rect -2238 -1775 -1426 -1774
rect -2238 -2575 -2237 -1775
rect -1427 -2575 -1426 -1775
rect 2172 -2573 2173 -1773
rect 2983 -2573 2984 -1773
rect 2172 -2574 2984 -2573
rect -2238 -2576 -1426 -2575
<< via4 >>
rect -2278 3144 -1416 3145
rect -2278 2295 -2277 3144
rect -2277 2295 -1417 3144
rect -1417 2295 -1416 3144
rect 2132 3144 2994 3145
rect 2132 2295 2133 3144
rect 2133 2295 2993 3144
rect 2993 2295 2994 3144
<< metal5 >>
rect -2302 3145 -1392 3169
rect -2302 2295 -2278 3145
rect -1416 2295 -1392 3145
rect 828 2683 1273 3152
rect 2108 3145 3018 3169
rect -2302 2271 -1392 2295
rect 2108 2295 2132 3145
rect 2994 2295 3018 3145
rect 2108 2271 3018 2295
use esd_diodes  esd_diodes_0
timestamp 1668294421
transform 1 0 -2972 0 -1 802
box 4520 -950 6580 2380
use esd_diodes  esd_diodes_1
timestamp 1668294421
transform 1 0 -7382 0 -1 802
box 4520 -950 6580 2380
use r_250  r_250_0
timestamp 1668438816
transform 1 0 53 0 1 53
box -53 -53 1220 3245
<< labels >>
rlabel metal2 165 2733 565 3133 6 in
port 1 n
rlabel metal1 -2272 1622 -1422 2289 0 vss
port 3 n
rlabel metal1 2138 1622 2988 2289 0 vss
rlabel metal1 -2232 -1770 -1432 -970 2 vdd
port 4 n
rlabel metal1 2178 -1768 2978 -968 6 vdd
rlabel metal5 828 2683 1273 3152 7 vss
rlabel metal2 168 182 565 579 7 out
port 2 n
<< end >>
