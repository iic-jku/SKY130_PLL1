magic
tech sky130A
magscale 1 2
timestamp 1666523630
<< error_p >>
rect 787 151 845 157
rect 787 117 799 151
rect 787 111 845 117
rect -845 -117 -787 -111
rect -845 -151 -833 -117
rect -845 -157 -787 -151
<< nwell >>
rect -1031 -289 1031 289
<< pmos >>
rect -831 -70 -801 70
rect -735 -70 -705 70
rect -639 -70 -609 70
rect -543 -70 -513 70
rect -447 -70 -417 70
rect -351 -70 -321 70
rect -255 -70 -225 70
rect -159 -70 -129 70
rect -63 -70 -33 70
rect 33 -70 63 70
rect 129 -70 159 70
rect 225 -70 255 70
rect 321 -70 351 70
rect 417 -70 447 70
rect 513 -70 543 70
rect 609 -70 639 70
rect 705 -70 735 70
rect 801 -70 831 70
<< pdiff >>
rect -893 58 -831 70
rect -893 -58 -881 58
rect -847 -58 -831 58
rect -893 -70 -831 -58
rect -801 58 -735 70
rect -801 -58 -785 58
rect -751 -58 -735 58
rect -801 -70 -735 -58
rect -705 58 -639 70
rect -705 -58 -689 58
rect -655 -58 -639 58
rect -705 -70 -639 -58
rect -609 58 -543 70
rect -609 -58 -593 58
rect -559 -58 -543 58
rect -609 -70 -543 -58
rect -513 58 -447 70
rect -513 -58 -497 58
rect -463 -58 -447 58
rect -513 -70 -447 -58
rect -417 58 -351 70
rect -417 -58 -401 58
rect -367 -58 -351 58
rect -417 -70 -351 -58
rect -321 58 -255 70
rect -321 -58 -305 58
rect -271 -58 -255 58
rect -321 -70 -255 -58
rect -225 58 -159 70
rect -225 -58 -209 58
rect -175 -58 -159 58
rect -225 -70 -159 -58
rect -129 58 -63 70
rect -129 -58 -113 58
rect -79 -58 -63 58
rect -129 -70 -63 -58
rect -33 58 33 70
rect -33 -58 -17 58
rect 17 -58 33 58
rect -33 -70 33 -58
rect 63 58 129 70
rect 63 -58 79 58
rect 113 -58 129 58
rect 63 -70 129 -58
rect 159 58 225 70
rect 159 -58 175 58
rect 209 -58 225 58
rect 159 -70 225 -58
rect 255 58 321 70
rect 255 -58 271 58
rect 305 -58 321 58
rect 255 -70 321 -58
rect 351 58 417 70
rect 351 -58 367 58
rect 401 -58 417 58
rect 351 -70 417 -58
rect 447 58 513 70
rect 447 -58 463 58
rect 497 -58 513 58
rect 447 -70 513 -58
rect 543 58 609 70
rect 543 -58 559 58
rect 593 -58 609 58
rect 543 -70 609 -58
rect 639 58 705 70
rect 639 -58 655 58
rect 689 -58 705 58
rect 639 -70 705 -58
rect 735 58 801 70
rect 735 -58 751 58
rect 785 -58 801 58
rect 735 -70 801 -58
rect 831 58 893 70
rect 831 -58 847 58
rect 881 -58 893 58
rect 831 -70 893 -58
<< pdiffc >>
rect -881 -58 -847 58
rect -785 -58 -751 58
rect -689 -58 -655 58
rect -593 -58 -559 58
rect -497 -58 -463 58
rect -401 -58 -367 58
rect -305 -58 -271 58
rect -209 -58 -175 58
rect -113 -58 -79 58
rect -17 -58 17 58
rect 79 -58 113 58
rect 175 -58 209 58
rect 271 -58 305 58
rect 367 -58 401 58
rect 463 -58 497 58
rect 559 -58 593 58
rect 655 -58 689 58
rect 751 -58 785 58
rect 847 -58 881 58
<< nsubdiff >>
rect -995 219 -899 253
rect 899 219 995 253
rect -995 157 -961 219
rect 961 157 995 219
rect -995 -219 -961 -157
rect 961 -219 995 -157
rect -995 -253 -899 -219
rect 899 -253 995 -219
<< nsubdiffcont >>
rect -899 219 899 253
rect -995 -157 -961 157
rect 961 -157 995 157
rect -899 -253 899 -219
<< poly >>
rect -753 151 -15 167
rect -753 117 -737 151
rect -703 117 -641 151
rect -607 117 -545 151
rect -511 117 -449 151
rect -415 117 -353 151
rect -319 117 -257 151
rect -223 117 -161 151
rect -127 117 -65 151
rect -31 117 -15 151
rect -753 101 -15 117
rect 399 151 561 167
rect 399 117 415 151
rect 449 117 511 151
rect 545 117 561 151
rect 399 101 561 117
rect 783 151 849 167
rect 783 117 799 151
rect 833 117 849 151
rect 783 101 849 117
rect -831 70 -801 96
rect -735 70 -705 101
rect -639 70 -609 101
rect -543 70 -513 101
rect -447 70 -417 101
rect -351 70 -321 101
rect -255 70 -225 101
rect -159 70 -129 101
rect -63 70 -33 101
rect 33 70 63 96
rect 129 70 159 96
rect 225 70 255 96
rect 321 70 351 96
rect 417 70 447 101
rect 513 70 543 101
rect 609 70 639 96
rect 705 70 735 96
rect 801 70 831 101
rect -831 -101 -801 -70
rect -735 -96 -705 -70
rect -639 -96 -609 -70
rect -543 -96 -513 -70
rect -447 -96 -417 -70
rect -351 -96 -321 -70
rect -255 -96 -225 -70
rect -159 -96 -129 -70
rect -63 -96 -33 -70
rect 33 -101 63 -70
rect 129 -101 159 -70
rect 225 -101 255 -70
rect 321 -101 351 -70
rect 417 -96 447 -70
rect 513 -96 543 -70
rect 609 -101 639 -70
rect 705 -101 735 -70
rect 801 -96 831 -70
rect -849 -117 -783 -101
rect -849 -151 -833 -117
rect -799 -151 -783 -117
rect -849 -167 -783 -151
rect 15 -117 369 -101
rect 15 -151 31 -117
rect 65 -151 127 -117
rect 161 -151 223 -117
rect 257 -151 319 -117
rect 353 -151 369 -117
rect 15 -167 369 -151
rect 591 -117 753 -101
rect 591 -151 607 -117
rect 641 -151 703 -117
rect 737 -151 753 -117
rect 591 -167 753 -151
<< polycont >>
rect -737 117 -703 151
rect -641 117 -607 151
rect -545 117 -511 151
rect -449 117 -415 151
rect -353 117 -319 151
rect -257 117 -223 151
rect -161 117 -127 151
rect -65 117 -31 151
rect 415 117 449 151
rect 511 117 545 151
rect 799 117 833 151
rect -833 -151 -799 -117
rect 31 -151 65 -117
rect 127 -151 161 -117
rect 223 -151 257 -117
rect 319 -151 353 -117
rect 607 -151 641 -117
rect 703 -151 737 -117
<< locali >>
rect -995 219 -899 253
rect 899 219 995 253
rect -995 157 -961 219
rect 961 157 995 219
rect -753 117 -737 151
rect -703 117 -641 151
rect -607 117 -545 151
rect -511 117 -449 151
rect -415 117 -353 151
rect -319 117 -257 151
rect -223 117 -161 151
rect -127 117 -65 151
rect -31 117 -15 151
rect 399 117 415 151
rect 449 117 511 151
rect 545 117 561 151
rect 783 117 799 151
rect 833 117 849 151
rect -881 58 -847 74
rect -881 -74 -847 -58
rect -785 58 -751 74
rect -785 -74 -751 -58
rect -689 58 -655 74
rect -689 -74 -655 -58
rect -593 58 -559 74
rect -593 -74 -559 -58
rect -497 58 -463 74
rect -497 -74 -463 -58
rect -401 58 -367 74
rect -401 -74 -367 -58
rect -305 58 -271 74
rect -305 -74 -271 -58
rect -209 58 -175 74
rect -209 -74 -175 -58
rect -113 58 -79 74
rect -113 -74 -79 -58
rect -17 58 17 74
rect -17 -74 17 -58
rect 79 58 113 74
rect 79 -74 113 -58
rect 175 58 209 74
rect 175 -74 209 -58
rect 271 58 305 74
rect 271 -74 305 -58
rect 367 58 401 74
rect 367 -74 401 -58
rect 463 58 497 74
rect 463 -74 497 -58
rect 559 58 593 74
rect 559 -74 593 -58
rect 655 58 689 74
rect 655 -74 689 -58
rect 751 58 785 74
rect 751 -74 785 -58
rect 847 58 881 74
rect 847 -74 881 -58
rect -849 -151 -833 -117
rect -799 -151 -783 -117
rect 15 -151 31 -117
rect 65 -151 127 -117
rect 161 -151 223 -117
rect 257 -151 319 -117
rect 353 -151 369 -117
rect 591 -151 607 -117
rect 641 -151 703 -117
rect 737 -151 753 -117
rect -995 -219 -961 -157
rect 961 -219 995 -157
rect -995 -253 -899 -219
rect 899 -253 995 -219
<< viali >>
rect -737 117 -703 151
rect -641 117 -607 151
rect -545 117 -511 151
rect -449 117 -415 151
rect -353 117 -319 151
rect -257 117 -223 151
rect -161 117 -127 151
rect -65 117 -31 151
rect 415 117 449 151
rect 511 117 545 151
rect 799 117 833 151
rect -881 -58 -847 58
rect -785 -58 -751 58
rect -689 -58 -655 58
rect -593 -58 -559 58
rect -497 -58 -463 58
rect -401 -58 -367 58
rect -305 -58 -271 58
rect -209 -58 -175 58
rect -113 -58 -79 58
rect -17 -58 17 58
rect 79 -58 113 58
rect 175 -58 209 58
rect 271 -58 305 58
rect 367 -58 401 58
rect 463 -58 497 58
rect 559 -58 593 58
rect 655 -58 689 58
rect 751 -58 785 58
rect 847 -58 881 58
rect -833 -151 -799 -117
rect 31 -151 65 -117
rect 127 -151 161 -117
rect 223 -151 257 -117
rect 319 -151 353 -117
rect 607 -151 641 -117
rect 703 -151 737 -117
<< metal1 >>
rect -749 151 -691 157
rect -653 151 -595 157
rect -557 151 -499 157
rect -461 151 -403 157
rect -365 151 -307 157
rect -269 151 -211 157
rect -173 151 -115 157
rect -77 151 -19 157
rect -749 117 -737 151
rect -703 117 -641 151
rect -607 117 -545 151
rect -511 117 -449 151
rect -415 117 -353 151
rect -319 117 -257 151
rect -223 117 -161 151
rect -127 117 -65 151
rect -31 117 -19 151
rect -749 111 -691 117
rect -653 111 -595 117
rect -557 111 -499 117
rect -461 111 -403 117
rect -365 111 -307 117
rect -269 111 -211 117
rect -173 111 -115 117
rect -77 111 -19 117
rect 403 151 461 157
rect 499 151 557 157
rect 403 117 415 151
rect 449 117 511 151
rect 545 117 557 151
rect 403 111 461 117
rect 499 111 557 117
rect 787 151 845 157
rect 787 117 799 151
rect 833 117 845 151
rect 787 111 845 117
rect -893 62 -739 70
rect -893 9 -890 62
rect -838 9 -794 62
rect -742 9 -739 62
rect -893 0 -881 9
rect -887 -58 -881 0
rect -847 0 -785 9
rect -847 -58 -841 0
rect -887 -70 -841 -58
rect -791 -58 -785 0
rect -751 0 -739 9
rect -695 58 -649 70
rect -695 0 -689 58
rect -751 -58 -745 0
rect -791 -70 -745 -58
rect -701 -9 -689 0
rect -655 0 -649 58
rect -605 62 -547 70
rect -605 9 -602 62
rect -550 9 -547 62
rect -605 0 -593 9
rect -655 -9 -643 0
rect -701 -62 -698 -9
rect -646 -62 -643 -9
rect -701 -70 -643 -62
rect -599 -58 -593 0
rect -559 0 -547 9
rect -503 58 -457 70
rect -503 0 -497 58
rect -559 -58 -553 0
rect -599 -70 -553 -58
rect -509 -9 -497 0
rect -463 0 -457 58
rect -413 62 -355 70
rect -413 9 -410 62
rect -358 9 -355 62
rect -413 0 -401 9
rect -463 -9 -451 0
rect -509 -62 -506 -9
rect -454 -62 -451 -9
rect -509 -70 -451 -62
rect -407 -58 -401 0
rect -367 0 -355 9
rect -311 58 -265 70
rect -311 0 -305 58
rect -367 -58 -361 0
rect -407 -70 -361 -58
rect -317 -9 -305 0
rect -271 0 -265 58
rect -221 62 -163 70
rect -221 9 -218 62
rect -166 9 -163 62
rect -221 0 -209 9
rect -271 -9 -259 0
rect -317 -62 -314 -9
rect -262 -62 -259 -9
rect -317 -70 -259 -62
rect -215 -58 -209 0
rect -175 0 -163 9
rect -119 58 -73 70
rect -119 0 -113 58
rect -175 -58 -169 0
rect -215 -70 -169 -58
rect -125 -9 -113 0
rect -79 0 -73 58
rect -29 62 29 70
rect -29 9 -26 62
rect 26 9 29 62
rect -29 0 -17 9
rect -79 -9 -67 0
rect -125 -62 -122 -9
rect -70 -62 -67 -9
rect -125 -70 -67 -62
rect -23 -58 -17 0
rect 17 0 29 9
rect 73 58 119 70
rect 73 0 79 58
rect 17 -58 23 0
rect -23 -70 23 -58
rect 67 -9 79 0
rect 113 0 119 58
rect 163 62 221 70
rect 163 9 166 62
rect 218 9 221 62
rect 163 0 175 9
rect 113 -9 125 0
rect 67 -62 70 -9
rect 122 -62 125 -9
rect 67 -70 125 -62
rect 169 -58 175 0
rect 209 0 221 9
rect 265 58 311 70
rect 265 0 271 58
rect 209 -58 215 0
rect 169 -70 215 -58
rect 259 -9 271 0
rect 305 0 311 58
rect 355 62 413 70
rect 355 9 358 62
rect 410 9 413 62
rect 355 0 367 9
rect 305 -9 317 0
rect 259 -62 262 -9
rect 314 -62 317 -9
rect 259 -70 317 -62
rect 361 -58 367 0
rect 401 0 413 9
rect 457 58 503 70
rect 457 0 463 58
rect 401 -58 407 0
rect 361 -70 407 -58
rect 451 -9 463 0
rect 497 0 503 58
rect 547 62 605 70
rect 547 9 550 62
rect 602 9 605 62
rect 547 0 559 9
rect 497 -9 509 0
rect 451 -62 454 -9
rect 506 -62 509 -9
rect 451 -70 509 -62
rect 553 -58 559 0
rect 593 0 605 9
rect 649 58 695 70
rect 649 0 655 58
rect 593 -58 599 0
rect 553 -70 599 -58
rect 643 -9 655 0
rect 689 0 695 58
rect 739 62 893 70
rect 739 9 742 62
rect 794 9 838 62
rect 890 9 893 62
rect 739 0 751 9
rect 689 -9 701 0
rect 643 -62 646 -9
rect 698 -62 701 -9
rect 643 -70 701 -62
rect 745 -58 751 0
rect 785 0 847 9
rect 785 -58 791 0
rect 745 -70 791 -58
rect 841 -58 847 0
rect 881 0 893 9
rect 881 -58 887 0
rect 841 -70 887 -58
rect -845 -117 -787 -111
rect -845 -151 -833 -117
rect -799 -151 -787 -117
rect -845 -157 -787 -151
rect 19 -117 77 -111
rect 115 -117 173 -111
rect 211 -117 269 -111
rect 307 -117 365 -111
rect 19 -151 31 -117
rect 65 -151 127 -117
rect 161 -151 223 -117
rect 257 -151 319 -117
rect 353 -151 365 -117
rect 19 -157 77 -151
rect 115 -157 173 -151
rect 211 -157 269 -151
rect 307 -157 365 -151
rect 595 -117 653 -111
rect 691 -117 749 -111
rect 595 -151 607 -117
rect 641 -151 703 -117
rect 737 -151 749 -117
rect 595 -157 653 -151
rect 691 -157 749 -151
<< via1 >>
rect -890 58 -838 62
rect -890 9 -881 58
rect -881 9 -847 58
rect -847 9 -838 58
rect -794 58 -742 62
rect -794 9 -785 58
rect -785 9 -751 58
rect -751 9 -742 58
rect -602 58 -550 62
rect -602 9 -593 58
rect -593 9 -559 58
rect -559 9 -550 58
rect -698 -58 -689 -9
rect -689 -58 -655 -9
rect -655 -58 -646 -9
rect -698 -62 -646 -58
rect -410 58 -358 62
rect -410 9 -401 58
rect -401 9 -367 58
rect -367 9 -358 58
rect -506 -58 -497 -9
rect -497 -58 -463 -9
rect -463 -58 -454 -9
rect -506 -62 -454 -58
rect -218 58 -166 62
rect -218 9 -209 58
rect -209 9 -175 58
rect -175 9 -166 58
rect -314 -58 -305 -9
rect -305 -58 -271 -9
rect -271 -58 -262 -9
rect -314 -62 -262 -58
rect -26 58 26 62
rect -26 9 -17 58
rect -17 9 17 58
rect 17 9 26 58
rect -122 -58 -113 -9
rect -113 -58 -79 -9
rect -79 -58 -70 -9
rect -122 -62 -70 -58
rect 166 58 218 62
rect 166 9 175 58
rect 175 9 209 58
rect 209 9 218 58
rect 70 -58 79 -9
rect 79 -58 113 -9
rect 113 -58 122 -9
rect 70 -62 122 -58
rect 358 58 410 62
rect 358 9 367 58
rect 367 9 401 58
rect 401 9 410 58
rect 262 -58 271 -9
rect 271 -58 305 -9
rect 305 -58 314 -9
rect 262 -62 314 -58
rect 550 58 602 62
rect 550 9 559 58
rect 559 9 593 58
rect 593 9 602 58
rect 454 -58 463 -9
rect 463 -58 497 -9
rect 497 -58 506 -9
rect 454 -62 506 -58
rect 742 58 794 62
rect 742 9 751 58
rect 751 9 785 58
rect 785 9 794 58
rect 838 58 890 62
rect 838 9 847 58
rect 847 9 881 58
rect 881 9 890 58
rect 646 -58 655 -9
rect 655 -58 689 -9
rect 689 -58 698 -9
rect 646 -62 698 -58
<< metal2 >>
rect -801 70 801 98
rect -893 62 893 70
rect -893 9 -890 62
rect -838 9 -794 62
rect -742 28 -602 62
rect -742 9 -739 28
rect -893 0 -739 9
rect -605 9 -602 28
rect -550 28 -410 62
rect -550 9 -547 28
rect -605 0 -547 9
rect -413 9 -410 28
rect -358 28 -218 62
rect -358 9 -355 28
rect -413 0 -355 9
rect -221 9 -218 28
rect -166 28 -26 62
rect -166 9 -163 28
rect -221 0 -163 9
rect -29 9 -26 28
rect 26 28 166 62
rect 26 9 29 28
rect -29 0 29 9
rect 163 9 166 28
rect 218 28 358 62
rect 218 9 221 28
rect 163 0 221 9
rect 355 9 358 28
rect 410 28 550 62
rect 410 9 413 28
rect 355 0 413 9
rect 547 9 550 28
rect 602 28 742 62
rect 602 9 605 28
rect 547 0 605 9
rect 739 9 742 28
rect 794 9 838 62
rect 890 9 893 62
rect 739 0 893 9
rect -701 -9 -643 0
rect -701 -62 -698 -9
rect -646 -28 -643 -9
rect -509 -9 -451 0
rect -509 -28 -506 -9
rect -646 -62 -506 -28
rect -454 -28 -451 -9
rect -317 -9 -259 0
rect -317 -28 -314 -9
rect -454 -62 -314 -28
rect -262 -28 -259 -9
rect -125 -9 -67 0
rect -125 -28 -122 -9
rect -262 -62 -122 -28
rect -70 -28 -67 -9
rect 67 -9 125 0
rect 67 -28 70 -9
rect -70 -62 70 -28
rect 122 -28 125 -9
rect 259 -9 317 0
rect 259 -28 262 -9
rect 122 -62 262 -28
rect 314 -28 317 -9
rect 451 -9 509 0
rect 451 -28 454 -9
rect 314 -62 454 -28
rect 506 -28 509 -9
rect 643 -9 701 0
rect 643 -28 646 -9
rect 506 -62 646 -28
rect 698 -62 701 -9
rect -701 -98 701 -62
<< properties >>
string FIXED_BBOX -978 -236 978 236
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.7 l 0.15 m 1 nf 18 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
