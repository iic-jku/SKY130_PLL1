magic
tech sky130A
magscale 1 2
timestamp 1668153059
<< metal1 >>
rect -1475 2104 6544 2304
rect -1475 1083 -1275 2104
rect -1105 1734 6174 1934
rect -1484 1074 -1266 1083
rect -1484 874 -1475 1074
rect -1275 874 -1266 1074
rect -1484 865 -1266 874
rect -1475 -3041 -1275 865
rect -1105 435 -905 1734
rect 5974 435 6174 1734
rect 6344 1083 6544 2104
rect 6335 1074 6553 1083
rect 6335 874 6344 1074
rect 6544 874 6553 1074
rect 6335 865 6553 874
rect -1114 426 -896 435
rect -1114 226 -1105 426
rect -905 226 -896 426
rect -1114 217 -896 226
rect 5965 426 6183 435
rect 5965 226 5974 426
rect 6174 226 6183 426
rect 5965 217 6183 226
rect -1105 -2393 -905 217
rect 2508 -135 2560 -129
rect 2508 -193 2560 -187
rect 2372 -416 2424 -410
rect 2372 -474 2424 -468
rect 2381 -1704 2415 -474
rect 2372 -1710 2424 -1704
rect 2372 -1768 2424 -1762
rect 2517 -1985 2551 -193
rect 2644 -518 2696 -512
rect 2644 -576 2696 -570
rect 2653 -1602 2687 -576
rect 2644 -1608 2696 -1602
rect 2644 -1666 2696 -1660
rect 2508 -1991 2560 -1985
rect 2508 -2049 2560 -2043
rect 5974 -2393 6174 217
rect -1114 -2402 -896 -2393
rect -1114 -2602 -1105 -2402
rect -905 -2602 -896 -2402
rect -1114 -2611 -896 -2602
rect 5965 -2402 6183 -2393
rect 5965 -2602 5974 -2402
rect 6174 -2602 6183 -2402
rect 5965 -2611 6183 -2602
rect -1484 -3050 -1266 -3041
rect -1484 -3250 -1475 -3050
rect -1275 -3250 -1266 -3050
rect -1484 -3259 -1266 -3250
rect -1475 -4282 -1275 -3259
rect -1105 -3912 -905 -2611
rect 5974 -3912 6174 -2611
rect 6344 -3041 6544 865
rect 6335 -3050 6553 -3041
rect 6335 -3250 6344 -3050
rect 6544 -3250 6553 -3050
rect 6335 -3259 6553 -3250
rect -1105 -4112 6174 -3912
rect 6344 -4282 6544 -3259
rect -1475 -4482 6544 -4282
<< via1 >>
rect -1475 874 -1275 1074
rect 6344 874 6544 1074
rect -1105 226 -905 426
rect 5974 226 6174 426
rect 2508 -187 2560 -135
rect 2372 -468 2424 -416
rect 2372 -1762 2424 -1710
rect 2644 -570 2696 -518
rect 2644 -1660 2696 -1608
rect 2508 -2043 2560 -1991
rect -1105 -2602 -905 -2402
rect 5974 -2602 6174 -2402
rect -1475 -3250 -1275 -3050
rect 6344 -3250 6544 -3050
<< metal2 >>
rect 1229 1295 1305 1305
rect 1229 1239 1239 1295
rect 1295 1239 1305 1295
rect 1229 1229 1305 1239
rect 2496 1293 2572 1303
rect 2496 1237 2506 1293
rect 2562 1282 2572 1293
rect 2562 1248 3818 1282
rect 2562 1237 2572 1248
rect 1250 1223 1284 1229
rect 2496 1227 2572 1237
rect 3784 1223 3818 1248
rect -1484 1074 -1266 1083
rect -1484 874 -1475 1074
rect -1275 874 -1266 1074
rect -1484 865 -1266 874
rect 6335 1074 6553 1083
rect 6335 874 6344 1074
rect 6544 874 6553 1074
rect 6335 865 6553 874
rect -1114 426 -896 435
rect -1114 226 -1105 426
rect -905 226 -896 426
rect -1114 217 -896 226
rect 5965 426 6183 435
rect 5965 226 5974 426
rect 6174 226 6183 426
rect 5965 217 6183 226
rect 1245 -37 1289 85
rect 2502 -187 2508 -135
rect 2560 -187 2566 -135
rect 2366 -468 2372 -416
rect 2424 -468 2430 -416
rect 2638 -570 2644 -518
rect 2696 -570 2702 -518
rect 2504 -1059 2564 -1050
rect 1228 -1119 1237 -1059
rect 1297 -1072 1306 -1059
rect 1297 -1106 2504 -1072
rect 1297 -1119 1306 -1106
rect 3762 -1072 3771 -1059
rect 2564 -1106 3771 -1072
rect 3762 -1119 3771 -1106
rect 3831 -1119 3840 -1059
rect 2504 -1128 2564 -1119
rect 2638 -1660 2644 -1608
rect 2696 -1660 2702 -1608
rect 2366 -1762 2372 -1710
rect 2424 -1762 2430 -1710
rect 2502 -2000 2508 -1991
rect 2484 -2034 2508 -2000
rect 2502 -2043 2508 -2034
rect 2560 -2000 2566 -1991
rect 2560 -2034 2586 -2000
rect 2560 -2043 2566 -2034
rect -1114 -2402 -896 -2393
rect -1114 -2602 -1105 -2402
rect -905 -2602 -896 -2402
rect -1114 -2611 -896 -2602
rect 5965 -2402 6183 -2393
rect 5965 -2602 5974 -2402
rect 6174 -2602 6183 -2402
rect 5965 -2611 6183 -2602
rect -1484 -3050 -1266 -3041
rect -1484 -3250 -1475 -3050
rect -1275 -3250 -1266 -3050
rect -1484 -3259 -1266 -3250
rect 6335 -3050 6553 -3041
rect 6335 -3250 6344 -3050
rect 6544 -3250 6553 -3050
rect 6335 -3259 6553 -3250
rect 1250 -3426 1284 -3401
rect 2496 -3415 2572 -3405
rect 3784 -3407 3818 -3401
rect 2496 -3426 2506 -3415
rect 1250 -3460 2506 -3426
rect 2496 -3471 2506 -3460
rect 2562 -3471 2572 -3415
rect 2496 -3481 2572 -3471
rect 3763 -3417 3839 -3407
rect 3763 -3473 3773 -3417
rect 3829 -3473 3839 -3417
rect 3763 -3483 3839 -3473
<< via2 >>
rect 1239 1239 1295 1295
rect 2506 1237 2562 1293
rect -1475 874 -1275 1074
rect 6344 874 6544 1074
rect -1105 226 -905 426
rect 5974 226 6174 426
rect 1237 -1119 1297 -1059
rect 2504 -1119 2564 -1059
rect 3771 -1119 3831 -1059
rect -1105 -2602 -905 -2402
rect 5974 -2602 6174 -2402
rect -1475 -3250 -1275 -3050
rect 6344 -3250 6544 -3050
rect 2506 -3471 2562 -3415
rect 3773 -3473 3829 -3417
<< metal3 >>
rect 1237 1311 1297 1342
rect 1223 1299 1311 1311
rect 1223 1235 1235 1299
rect 1299 1235 1311 1299
rect 1223 1223 1311 1235
rect 2490 1297 2578 1309
rect 2490 1233 2502 1297
rect 2566 1294 2578 1297
rect 2566 1234 2609 1294
rect 2566 1233 2578 1234
rect 2490 1221 2578 1233
rect -1484 1074 -1266 1083
rect -1484 874 -1475 1074
rect -1275 1003 -1266 1074
rect 6335 1074 6553 1083
rect 6335 1003 6344 1074
rect -1275 943 -716 1003
rect 5784 943 6344 1003
rect -1275 874 -1266 943
rect -1484 865 -1266 874
rect 6335 874 6344 943
rect 6544 874 6553 1074
rect 6335 865 6553 874
rect -1114 426 -896 435
rect -1114 226 -1105 426
rect -905 355 -896 426
rect 5965 426 6183 435
rect 5965 355 5974 426
rect -905 295 -716 355
rect 5784 295 5974 355
rect -905 226 -896 295
rect -1114 217 -896 226
rect 5965 226 5974 295
rect 6174 226 6183 426
rect 5965 217 6183 226
rect 1223 73 1311 85
rect 1223 9 1235 73
rect 1299 9 1311 73
rect 1223 -3 1311 9
rect 2490 73 2578 85
rect 2490 9 2502 73
rect 2566 9 2578 73
rect 2490 -3 2578 9
rect 537 -140 597 -107
rect 528 -147 606 -140
rect 528 -211 535 -147
rect 599 -211 606 -147
rect 528 -218 606 -211
rect 537 -1046 597 -218
rect 537 -1180 597 -1132
rect 528 -1187 606 -1180
rect 528 -1251 535 -1187
rect 599 -1251 606 -1187
rect 528 -1258 606 -1251
rect 537 -2071 597 -1258
rect 834 -1440 894 -107
rect 1237 -1054 1297 -3
rect 1232 -1059 1302 -1054
rect 1232 -1119 1237 -1059
rect 1297 -1119 1302 -1059
rect 1232 -1124 1302 -1119
rect 1639 -1180 1699 -107
rect 1936 -400 1996 -107
rect 1927 -407 2005 -400
rect 1927 -471 1934 -407
rect 1998 -471 2005 -407
rect 1927 -478 2005 -471
rect 1936 -1046 1996 -478
rect 2504 -1054 2564 -3
rect 3072 -660 3132 -107
rect 3369 -140 3429 -107
rect 3360 -147 3438 -140
rect 3360 -211 3367 -147
rect 3431 -211 3438 -147
rect 3360 -218 3438 -211
rect 3369 -600 3429 -218
rect 4174 -400 4234 -107
rect 4165 -407 4243 -400
rect 4165 -471 4172 -407
rect 4236 -471 4243 -407
rect 4165 -478 4243 -471
rect 3063 -667 3141 -660
rect 3063 -731 3070 -667
rect 3134 -731 3141 -667
rect 3063 -738 3141 -731
rect 3360 -667 3438 -660
rect 3360 -731 3367 -667
rect 3431 -731 3438 -667
rect 3360 -738 3438 -731
rect 3072 -1046 3132 -738
rect 2499 -1059 2569 -1054
rect 2499 -1119 2504 -1059
rect 2564 -1119 2569 -1059
rect 2499 -1124 2569 -1119
rect 1630 -1187 1708 -1180
rect 1630 -1251 1637 -1187
rect 1701 -1251 1708 -1187
rect 1630 -1258 1708 -1251
rect 825 -1447 903 -1440
rect 825 -1511 832 -1447
rect 896 -1511 903 -1447
rect 825 -1518 903 -1511
rect 834 -1960 894 -1578
rect 1639 -1700 1699 -1318
rect 1936 -1440 1996 -1132
rect 1927 -1447 2005 -1440
rect 1927 -1511 1934 -1447
rect 1998 -1511 2005 -1447
rect 1927 -1518 2005 -1511
rect 1630 -1707 1708 -1700
rect 1630 -1771 1637 -1707
rect 1701 -1771 1708 -1707
rect 1630 -1778 1708 -1771
rect 825 -1967 903 -1960
rect 825 -2031 832 -1967
rect 896 -2031 903 -1967
rect 825 -2038 903 -2031
rect 834 -2071 894 -2038
rect 1639 -2071 1699 -1778
rect 1936 -2071 1996 -1518
rect 2504 -2175 2564 -1124
rect 3072 -1960 3132 -1132
rect 3063 -1967 3141 -1960
rect 3063 -2031 3070 -1967
rect 3134 -2031 3141 -1967
rect 3063 -2038 3141 -2031
rect 3072 -2071 3132 -2038
rect 3369 -2071 3429 -738
rect 4174 -860 4234 -478
rect 4471 -920 4531 -107
rect 4165 -927 4243 -920
rect 4165 -991 4172 -927
rect 4236 -991 4243 -927
rect 4165 -998 4243 -991
rect 4462 -927 4540 -920
rect 4462 -991 4469 -927
rect 4533 -991 4540 -927
rect 4462 -998 4540 -991
rect 3766 -1059 3836 -1054
rect 3766 -1119 3771 -1059
rect 3831 -1119 3836 -1059
rect 3766 -1124 3836 -1119
rect 3771 -2175 3831 -1124
rect 4174 -2071 4234 -998
rect 4471 -1046 4531 -998
rect 4471 -1700 4531 -1132
rect 4462 -1707 4540 -1700
rect 4462 -1771 4469 -1707
rect 4533 -1771 4540 -1707
rect 4462 -1778 4540 -1771
rect 4471 -2071 4531 -1778
rect 2490 -2187 2578 -2175
rect 2490 -2251 2502 -2187
rect 2566 -2251 2578 -2187
rect 2490 -2263 2578 -2251
rect 3757 -2187 3845 -2175
rect 3757 -2251 3769 -2187
rect 3833 -2251 3845 -2187
rect 3757 -2263 3845 -2251
rect -1114 -2402 -896 -2393
rect -1114 -2602 -1105 -2402
rect -905 -2473 -896 -2402
rect 5965 -2402 6183 -2393
rect 5965 -2473 5974 -2402
rect -905 -2533 -716 -2473
rect 5784 -2533 5974 -2473
rect -905 -2602 -896 -2533
rect -1114 -2611 -896 -2602
rect 5965 -2602 5974 -2533
rect 6174 -2602 6183 -2402
rect 5965 -2611 6183 -2602
rect -1484 -3050 -1266 -3041
rect -1484 -3250 -1475 -3050
rect -1275 -3121 -1266 -3050
rect 6335 -3050 6553 -3041
rect 6335 -3121 6344 -3050
rect -1275 -3181 -716 -3121
rect 5784 -3181 6344 -3121
rect -1275 -3250 -1266 -3181
rect -1484 -3259 -1266 -3250
rect 6335 -3250 6344 -3181
rect 6544 -3250 6553 -3050
rect 6335 -3259 6553 -3250
rect 2490 -3411 2578 -3399
rect 2490 -3412 2502 -3411
rect 2459 -3472 2502 -3412
rect 2490 -3475 2502 -3472
rect 2566 -3475 2578 -3411
rect 2490 -3487 2578 -3475
rect 3757 -3413 3845 -3401
rect 3757 -3477 3769 -3413
rect 3833 -3477 3845 -3413
rect 3757 -3489 3845 -3477
rect 3771 -3520 3831 -3489
<< via3 >>
rect 1235 1295 1299 1299
rect 1235 1239 1239 1295
rect 1239 1239 1295 1295
rect 1295 1239 1299 1295
rect 1235 1235 1299 1239
rect 2502 1293 2566 1297
rect 2502 1237 2506 1293
rect 2506 1237 2562 1293
rect 2562 1237 2566 1293
rect 2502 1233 2566 1237
rect 1235 9 1299 73
rect 2502 9 2566 73
rect 535 -211 599 -147
rect 535 -1251 599 -1187
rect 1934 -471 1998 -407
rect 3367 -211 3431 -147
rect 4172 -471 4236 -407
rect 3070 -731 3134 -667
rect 3367 -731 3431 -667
rect 1637 -1251 1701 -1187
rect 832 -1511 896 -1447
rect 1934 -1511 1998 -1447
rect 1637 -1771 1701 -1707
rect 832 -2031 896 -1967
rect 3070 -2031 3134 -1967
rect 4172 -991 4236 -927
rect 4469 -991 4533 -927
rect 4469 -1771 4533 -1707
rect 2502 -2251 2566 -2187
rect 3769 -2251 3833 -2187
rect 2502 -3415 2566 -3411
rect 2502 -3471 2506 -3415
rect 2506 -3471 2562 -3415
rect 2562 -3471 2566 -3415
rect 2502 -3475 2566 -3471
rect 3769 -3417 3833 -3413
rect 3769 -3473 3773 -3417
rect 3773 -3473 3829 -3417
rect 3829 -3473 3833 -3417
rect 3769 -3477 3833 -3473
<< metal4 >>
rect 1223 1299 1311 1311
rect 686 1221 746 1281
rect 1223 1235 1235 1299
rect 1299 1235 1311 1299
rect 2490 1297 2578 1309
rect 1223 1223 1311 1235
rect 1237 85 1297 1223
rect 1788 1221 1848 1281
rect 2490 1233 2502 1297
rect 2566 1233 2578 1297
rect 2490 1221 2578 1233
rect 3220 1221 3280 1281
rect 4322 1221 4382 1281
rect 2504 85 2564 1221
rect 1223 73 1311 85
rect 1223 9 1235 73
rect 1299 9 1311 73
rect 1223 -3 1311 9
rect 2490 73 2578 85
rect 2490 9 2502 73
rect 2566 9 2578 73
rect 2490 -3 2578 9
rect 528 -147 606 -140
rect 528 -149 535 -147
rect 0 -209 535 -149
rect 528 -211 535 -209
rect 599 -149 606 -147
rect 3360 -147 3438 -140
rect 3360 -149 3367 -147
rect 599 -209 3367 -149
rect 599 -211 606 -209
rect 528 -218 606 -211
rect 3360 -211 3367 -209
rect 3431 -149 3438 -147
rect 3431 -209 5068 -149
rect 3431 -211 3438 -209
rect 3360 -218 3438 -211
rect 1927 -407 2005 -400
rect 1927 -409 1934 -407
rect 0 -469 1934 -409
rect 1927 -471 1934 -469
rect 1998 -409 2005 -407
rect 4165 -407 4243 -400
rect 4165 -409 4172 -407
rect 1998 -469 4172 -409
rect 1998 -471 2005 -469
rect 1927 -478 2005 -471
rect 4165 -471 4172 -469
rect 4236 -409 4243 -407
rect 4236 -469 5068 -409
rect 4236 -471 4243 -469
rect 4165 -478 4243 -471
rect 3063 -667 3141 -660
rect 3063 -669 3070 -667
rect 0 -729 3070 -669
rect 3063 -731 3070 -729
rect 3134 -669 3141 -667
rect 3360 -667 3438 -660
rect 3360 -669 3367 -667
rect 3134 -729 3367 -669
rect 3134 -731 3141 -729
rect 3063 -738 3141 -731
rect 3360 -731 3367 -729
rect 3431 -669 3438 -667
rect 3431 -729 5068 -669
rect 3431 -731 3438 -729
rect 3360 -738 3438 -731
rect 4165 -927 4243 -920
rect 4165 -929 4172 -927
rect 0 -989 4172 -929
rect 4165 -991 4172 -989
rect 4236 -929 4243 -927
rect 4462 -927 4540 -920
rect 4462 -929 4469 -927
rect 4236 -989 4469 -929
rect 4236 -991 4243 -989
rect 4165 -998 4243 -991
rect 4462 -991 4469 -989
rect 4533 -929 4540 -927
rect 4533 -989 5068 -929
rect 4533 -991 4540 -989
rect 4462 -998 4540 -991
rect 528 -1187 606 -1180
rect 528 -1189 535 -1187
rect 0 -1249 535 -1189
rect 528 -1251 535 -1249
rect 599 -1189 606 -1187
rect 1630 -1187 1708 -1180
rect 1630 -1189 1637 -1187
rect 599 -1249 1637 -1189
rect 599 -1251 606 -1249
rect 528 -1258 606 -1251
rect 1630 -1251 1637 -1249
rect 1701 -1189 1708 -1187
rect 1701 -1249 5068 -1189
rect 1701 -1251 1708 -1249
rect 1630 -1258 1708 -1251
rect 825 -1447 903 -1440
rect 825 -1449 832 -1447
rect 0 -1509 832 -1449
rect 825 -1511 832 -1509
rect 896 -1449 903 -1447
rect 1927 -1447 2005 -1440
rect 1927 -1449 1934 -1447
rect 896 -1509 1934 -1449
rect 896 -1511 903 -1509
rect 825 -1518 903 -1511
rect 1927 -1511 1934 -1509
rect 1998 -1449 2005 -1447
rect 1998 -1509 5068 -1449
rect 1998 -1511 2005 -1509
rect 1927 -1518 2005 -1511
rect 1630 -1707 1708 -1700
rect 1630 -1709 1637 -1707
rect 0 -1769 1637 -1709
rect 1630 -1771 1637 -1769
rect 1701 -1709 1708 -1707
rect 4462 -1707 4540 -1700
rect 4462 -1709 4469 -1707
rect 1701 -1769 4469 -1709
rect 1701 -1771 1708 -1769
rect 1630 -1778 1708 -1771
rect 4462 -1771 4469 -1769
rect 4533 -1709 4540 -1707
rect 4533 -1769 5068 -1709
rect 4533 -1771 4540 -1769
rect 4462 -1778 4540 -1771
rect 825 -1967 903 -1960
rect 825 -1969 832 -1967
rect 0 -2029 832 -1969
rect 825 -2031 832 -2029
rect 896 -1969 903 -1967
rect 3063 -1967 3141 -1960
rect 3063 -1969 3070 -1967
rect 896 -2029 3070 -1969
rect 896 -2031 903 -2029
rect 825 -2038 903 -2031
rect 3063 -2031 3070 -2029
rect 3134 -1969 3141 -1967
rect 3134 -2029 5068 -1969
rect 3134 -2031 3141 -2029
rect 3063 -2038 3141 -2031
rect 2490 -2187 2578 -2175
rect 2490 -2251 2502 -2187
rect 2566 -2251 2578 -2187
rect 2490 -2263 2578 -2251
rect 3757 -2187 3845 -2175
rect 3757 -2251 3769 -2187
rect 3833 -2251 3845 -2187
rect 3757 -2263 3845 -2251
rect 2504 -3399 2564 -2263
rect 686 -3459 746 -3399
rect 1788 -3459 1848 -3399
rect 2490 -3411 2578 -3399
rect 2490 -3475 2502 -3411
rect 2566 -3475 2578 -3411
rect 3220 -3459 3280 -3399
rect 3771 -3401 3831 -2263
rect 3757 -3413 3845 -3401
rect 2490 -3487 2578 -3475
rect 3757 -3477 3769 -3413
rect 3833 -3477 3845 -3413
rect 4322 -3459 4382 -3399
rect 3757 -3489 3845 -3477
use delay_cell_4  delay_cell_4_0
timestamp 1668153059
transform 1 0 865 0 1 138
box -1581 -735 1669 1085
use delay_cell_4  delay_cell_4_1
timestamp 1668153059
transform -1 0 4203 0 1 138
box -1581 -735 1669 1085
use delay_cell_4  delay_cell_4_2
timestamp 1668153059
transform -1 0 4203 0 -1 -2316
box -1581 -735 1669 1085
use delay_cell_4  delay_cell_4_3
timestamp 1668153059
transform 1 0 865 0 -1 -2316
box -1581 -735 1669 1085
<< labels >>
rlabel metal4 686 1221 746 1281 0 inv1
rlabel metal4 1788 1221 1848 1281 0 inv2
rlabel metal4 3220 1221 3280 1281 0 inv3
rlabel metal4 4322 1221 4382 1281 6 inv4
rlabel metal4 528 -218 606 -140 0 out1
port 6 n
rlabel metal4 1927 -478 2005 -400 0 out2
port 7 n
rlabel metal4 3063 -738 3141 -660 7 out3
port 8 n
rlabel metal4 4462 -998 4540 -920 0 out4
port 9 n
rlabel metal4 528 -1258 606 -1180 0 out8
port 13 n
rlabel metal1 2653 -1106 2687 -1072 7 b2
port 3 n
rlabel metal1 2517 -1106 2551 -1072 0 b1
port 4 n
rlabel metal1 2381 -1106 2415 -1072 0 b0
port 5 n
rlabel metal4 1927 -1518 2005 -1440 5 out7
port 12 n
rlabel metal4 4462 -1778 4540 -1700 0 out5
port 10 n
rlabel metal4 3063 -2038 3141 -1960 3 out6
port 11 n
rlabel metal4 4322 -3459 4382 -3399 7 inv5
rlabel metal4 3220 -3459 3280 -3399 3 inv6
rlabel metal4 1788 -3459 1848 -3399 4 inv7
rlabel metal4 686 -3459 746 -3399 7 inv8
rlabel metal3 5784 943 5844 1003 0 vdd
port 1 n
rlabel metal3 5784 -3181 5844 -3121 0 vdd
rlabel metal3 5784 295 5844 355 0 vss
port 2 n
rlabel metal3 5784 -2533 5844 -2473 0 vss
rlabel metal3 -776 943 -716 1003 7 vdd
rlabel metal3 -776 295 -716 355 0 vss
rlabel metal3 -776 -2533 -716 -2473 0 vss
rlabel metal3 -776 -3181 -716 -3121 3 vdd
rlabel metal2 1362 -1106 1396 -1072 0 vdelay
port 14 n
<< end >>
