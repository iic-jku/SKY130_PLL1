magic
tech sky130A
magscale 1 2
timestamp 1652803914
<< nwell >>
rect -228 -53 -53 525
<< metal1 >>
rect -217 396 -153 402
rect -217 387 -211 396
rect -228 353 -211 387
rect -217 344 -211 353
rect -159 387 -153 396
rect -159 353 -53 387
rect -159 344 -153 353
rect -217 338 -153 344
rect -228 85 -102 119
rect -136 -89 -102 85
rect 148 -80 212 -74
rect 148 -89 154 -80
rect -136 -123 154 -89
rect 148 -132 154 -123
rect 206 -132 212 -80
rect 148 -138 212 -132
rect -125 -432 -61 -426
rect -125 -441 -119 -432
rect -324 -475 -119 -441
rect -125 -484 -119 -475
rect -67 -441 -61 -432
rect -67 -475 -53 -441
rect -67 -484 -61 -475
rect -125 -490 -61 -484
<< via1 >>
rect -211 344 -159 396
rect 154 -132 206 -80
rect -119 -484 -67 -432
<< metal2 >>
rect -217 396 -153 402
rect -217 344 -211 396
rect -159 344 -153 396
rect -217 338 -153 344
rect -946 -123 -681 -89
rect -202 -336 -168 338
rect -130 304 -56 313
rect -130 248 -121 304
rect -65 248 -56 304
rect -130 239 -56 248
rect -222 -345 -148 -336
rect -222 -401 -213 -345
rect -157 -401 -148 -345
rect -222 -410 -148 -401
rect -110 -426 -76 239
rect 148 -80 212 -74
rect 148 -132 154 -80
rect 206 -132 212 -80
rect 148 -138 212 -132
rect -125 -432 -61 -426
rect -125 -484 -119 -432
rect -67 -484 -61 -432
rect -125 -490 -61 -484
<< via2 >>
rect -121 248 -65 304
rect -213 -401 -157 -345
<< metal3 >>
rect -130 306 -56 313
rect -228 304 -53 306
rect -228 248 -121 304
rect -65 248 -53 304
rect -228 246 -53 248
rect -130 239 -56 246
rect -222 -343 -148 -336
rect -324 -345 -53 -343
rect -324 -401 -213 -345
rect -157 -401 -53 -345
rect -324 -403 -53 -401
rect -222 -410 -148 -403
use n_buf  sky130_fd_pr__nfet_01v8_5ZA63U_0
timestamp 1652802656
transform 1 0 258 0 1 -333
box -311 -280 311 280
use n_buf  sky130_fd_pr__nfet_01v8_5ZA63U_1
timestamp 1652802656
transform 1 0 -635 0 1 -333
box -311 -280 311 280
use p_buf  sky130_fd_pr__pfet_01v8_X679XQ_0
timestamp 1652802024
transform 1 0 306 0 1 236
box -359 -289 359 289
use p_buf  sky130_fd_pr__pfet_01v8_X679XQ_1
timestamp 1652802024
transform 1 0 -587 0 1 236
box -359 -289 359 289
<< end >>
