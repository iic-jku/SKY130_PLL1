magic
tech sky130A
magscale 1 2
timestamp 1668357910
<< pwell >>
rect -359 -280 359 280
<< nmos >>
rect -159 -70 -129 70
rect -63 -70 -33 70
rect 33 -70 63 70
rect 129 -70 159 70
<< ndiff >>
rect -221 58 -159 70
rect -221 -58 -209 58
rect -175 -58 -159 58
rect -221 -70 -159 -58
rect -129 58 -63 70
rect -129 -58 -113 58
rect -79 -58 -63 58
rect -129 -70 -63 -58
rect -33 58 33 70
rect -33 -58 -17 58
rect 17 -58 33 58
rect -33 -70 33 -58
rect 63 58 129 70
rect 63 -58 79 58
rect 113 -58 129 58
rect 63 -70 129 -58
rect 159 58 221 70
rect 159 -58 175 58
rect 209 -58 221 58
rect 159 -70 221 -58
<< ndiffc >>
rect -209 -58 -175 58
rect -113 -58 -79 58
rect -17 -58 17 58
rect 79 -58 113 58
rect 175 -58 209 58
<< psubdiff >>
rect -323 210 -227 244
rect 227 210 323 244
rect -323 148 -289 210
rect 289 148 323 210
rect -323 -210 -289 -148
rect 289 -210 323 -148
rect -323 -244 -227 -210
rect 227 -244 323 -210
<< psubdiffcont >>
rect -227 210 227 244
rect -323 -148 -289 148
rect 289 -148 323 148
rect -227 -244 227 -210
<< poly >>
rect -81 142 81 158
rect -81 108 -65 142
rect -31 108 31 142
rect 65 108 81 142
rect -159 70 -129 96
rect -81 92 81 108
rect -63 70 -33 92
rect 33 70 63 92
rect 129 70 159 96
rect -159 -92 -129 -70
rect -177 -108 -111 -92
rect -63 -96 -33 -70
rect 33 -96 63 -70
rect 129 -92 159 -70
rect -177 -142 -161 -108
rect -127 -142 -111 -108
rect -177 -158 -111 -142
rect 111 -108 177 -92
rect 111 -142 127 -108
rect 161 -142 177 -108
rect 111 -158 177 -142
<< polycont >>
rect -65 108 -31 142
rect 31 108 65 142
rect -161 -142 -127 -108
rect 127 -142 161 -108
<< locali >>
rect -323 210 -227 244
rect 227 210 323 244
rect -323 148 -289 210
rect 289 148 323 210
rect -81 108 -65 142
rect -31 108 31 142
rect 65 108 81 142
rect -209 58 -175 74
rect -209 -74 -175 -58
rect -113 58 -79 74
rect -113 -74 -79 -58
rect -17 58 17 74
rect -17 -74 17 -58
rect 79 58 113 74
rect 79 -74 113 -58
rect 175 58 209 74
rect 175 -74 209 -58
rect -177 -142 -161 -108
rect -127 -142 -111 -108
rect 111 -142 127 -108
rect 161 -142 177 -108
rect -323 -210 -289 -148
rect 289 -210 323 -148
rect -323 -244 -227 -210
rect 227 -244 323 -210
<< viali >>
rect -65 108 -31 142
rect 31 108 65 142
rect -209 -58 -175 58
rect -113 -58 -79 58
rect -17 -58 17 58
rect 79 -58 113 58
rect 175 -58 209 58
rect -161 -142 -127 -108
rect 127 -142 161 -108
<< metal1 >>
rect -77 142 -19 148
rect 19 142 77 148
rect -81 108 -65 142
rect -31 108 31 142
rect 65 108 81 142
rect -77 102 -19 108
rect 19 102 77 108
rect -215 58 -169 70
rect -215 0 -209 58
rect -221 -8 -209 0
rect -175 0 -169 58
rect -119 58 -73 70
rect -119 0 -113 58
rect -175 -8 -113 0
rect -79 0 -73 58
rect -29 61 29 70
rect -29 8 -26 61
rect 26 8 29 61
rect -29 0 -17 8
rect -79 -8 -67 0
rect -221 -61 -218 -8
rect -166 -61 -122 -8
rect -70 -61 -67 -8
rect -221 -70 -67 -61
rect -23 -58 -17 0
rect 17 0 29 8
rect 73 58 119 70
rect 73 0 79 58
rect 17 -58 23 0
rect -23 -70 23 -58
rect 67 -8 79 0
rect 113 0 119 58
rect 169 58 215 70
rect 169 0 175 58
rect 113 -8 175 0
rect 209 0 215 58
rect 209 -8 221 0
rect 67 -61 70 -8
rect 122 -61 166 -8
rect 218 -61 221 -8
rect 67 -70 221 -61
rect -210 -102 -173 -70
rect 172 -102 209 -70
rect -210 -108 -115 -102
rect -210 -142 -161 -108
rect -127 -142 -115 -108
rect -210 -148 -115 -142
rect 115 -108 209 -102
rect 115 -142 127 -108
rect 161 -142 209 -108
rect 115 -148 209 -142
<< via1 >>
rect -26 58 26 61
rect -26 8 -17 58
rect -17 8 17 58
rect 17 8 26 58
rect -218 -58 -209 -8
rect -209 -58 -175 -8
rect -175 -58 -166 -8
rect -218 -61 -166 -58
rect -122 -58 -113 -8
rect -113 -58 -79 -8
rect -79 -58 -70 -8
rect -122 -61 -70 -58
rect 70 -58 79 -8
rect 79 -58 113 -8
rect 113 -58 122 -8
rect 70 -61 122 -58
rect 166 -58 175 -8
rect 175 -58 209 -8
rect 209 -58 218 -8
rect 166 -61 218 -58
<< metal2 >>
rect -29 61 29 70
rect -29 8 -26 61
rect 26 8 29 61
rect -29 0 29 8
rect -221 -8 -67 0
rect -221 -61 -218 -8
rect -166 -61 -122 -8
rect -70 -28 -67 -8
rect 67 -8 221 0
rect 67 -28 70 -8
rect -70 -61 70 -28
rect 122 -61 166 -8
rect 218 -61 221 -8
rect -221 -70 221 -61
<< properties >>
string FIXED_BBOX -306 -227 306 227
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.7 l 0.150 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
