magic
tech sky130A
magscale 1 2
timestamp 1668153059
<< metal3 >>
rect 0 64100 100 70200
rect 6600 64100 6700 70200
rect 13200 64100 13300 70200
rect 19800 64100 19900 70200
rect 26400 64100 26500 70200
rect 33000 64100 33100 70200
rect 39600 64100 39700 70200
rect 46200 64100 46300 70200
rect 52800 64100 52900 70200
rect 59400 64100 59500 70200
rect 0 64000 65599 64100
rect 0 57700 100 64000
rect 6600 57700 6700 64000
rect 13200 57700 13300 64000
rect 19800 57700 19900 64000
rect 26400 57700 26500 64000
rect 33000 57700 33100 64000
rect 39600 57700 39700 64000
rect 46200 57700 46300 64000
rect 52800 57700 52900 64000
rect 59400 57700 59500 64000
rect 0 57600 65599 57700
rect 0 51300 100 57600
rect 6600 51300 6700 57600
rect 13200 51300 13300 57600
rect 19800 51300 19900 57600
rect 26400 51300 26500 57600
rect 33000 51300 33100 57600
rect 39600 51300 39700 57600
rect 46200 51300 46300 57600
rect 52800 51300 52900 57600
rect 59400 51300 59500 57600
rect 0 51200 65599 51300
rect 0 44900 100 51200
rect 6600 44900 6700 51200
rect 13200 44900 13300 51200
rect 19800 44900 19900 51200
rect 26400 44900 26500 51200
rect 33000 44900 33100 51200
rect 39600 44900 39700 51200
rect 46200 44900 46300 51200
rect 52800 44900 52900 51200
rect 59400 44900 59500 51200
rect 0 44800 65599 44900
rect 0 38500 100 44800
rect 6600 38500 6700 44800
rect 13200 38500 13300 44800
rect 19800 38500 19900 44800
rect 26400 38500 26500 44800
rect 33000 38500 33100 44800
rect 39600 38500 39700 44800
rect 46200 38500 46300 44800
rect 52800 38500 52900 44800
rect 59400 38500 59500 44800
rect 0 38400 65599 38500
rect 0 32100 100 38400
rect 6600 32100 6700 38400
rect 13200 32100 13300 38400
rect 19800 32100 19900 38400
rect 26400 32100 26500 38400
rect 33000 32100 33100 38400
rect 39600 32100 39700 38400
rect 46200 32100 46300 38400
rect 52800 32100 52900 38400
rect 59400 32100 59500 38400
rect 0 32000 65599 32100
rect 0 25700 100 32000
rect 6600 25700 6700 32000
rect 13200 25700 13300 32000
rect 19800 25700 19900 32000
rect 26400 25700 26500 32000
rect 33000 25700 33100 32000
rect 39600 25700 39700 32000
rect 46200 25700 46300 32000
rect 52800 25700 52900 32000
rect 59400 25700 59500 32000
rect 0 25600 65599 25700
rect 0 19300 100 25600
rect 6600 19300 6700 25600
rect 13200 19300 13300 25600
rect 19800 19300 19900 25600
rect 26400 19300 26500 25600
rect 33000 19300 33100 25600
rect 39600 19300 39700 25600
rect 46200 19300 46300 25600
rect 52800 19300 52900 25600
rect 59400 19300 59500 25600
rect 0 19200 65599 19300
rect 0 12900 100 19200
rect 6600 12900 6700 19200
rect 13200 12900 13300 19200
rect 19800 12900 19900 19200
rect 26400 12900 26500 19200
rect 33000 12900 33100 19200
rect 39600 12900 39700 19200
rect 46200 12900 46300 19200
rect 52800 12900 52900 19200
rect 59400 12900 59500 19200
rect 0 12800 65599 12900
rect 0 6500 100 12800
rect 6600 6500 6700 12800
rect 13200 6500 13300 12800
rect 19800 6500 19900 12800
rect 26400 6500 26500 12800
rect 33000 6500 33100 12800
rect 39600 6500 39700 12800
rect 46200 6500 46300 12800
rect 52800 6500 52900 12800
rect 59400 6500 59500 12800
rect 0 6400 65599 6500
rect 0 100 100 6400
rect 6600 100 6700 6400
rect 13200 100 13300 6400
rect 19800 100 19900 6400
rect 26400 100 26500 6400
rect 33000 100 33100 6400
rect 39600 100 39700 6400
rect 46200 100 46300 6400
rect 52800 100 52900 6400
rect 59400 100 59500 6400
rect 0 0 65599 100
<< metal4 >>
rect -96 70200 65695 70296
rect -96 0 0 70200
rect 6199 0 6295 70200
rect 12799 0 12895 70200
rect 19399 0 19495 70200
rect 25999 0 26095 70200
rect 32599 0 32695 70200
rect 39199 0 39295 70200
rect 45799 0 45895 70200
rect 52399 70088 52498 70200
rect 52402 111 52498 70088
rect 52399 0 52498 111
rect 58999 0 59095 70200
rect 65599 0 65695 70200
rect -96 -96 65695 0
use sky130_fd_pr__cap_mim_m3_1_LJ5JLG  sky130_fd_pr__cap_mim_m3_1_LJ5JLG_0
array 0 9 6600 0 10 6400
timestamp 1668153059
transform 1 0 3150 0 1 3100
box -3150 -3100 3149 3100
<< end >>
