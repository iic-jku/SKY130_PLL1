* SPICE3 file created from core_complete_1.ext - technology: sky130A
V1 vdd vss 1.8
V2 vb1 vss 0.6
V3 vb2 vss 0.6
V4 vss gnd 0
V10 bit0 vss 1.8 
*ss
V11 bit1 vss 0 
*tt
V12 bit2 vss 1.8 
*ff

.subckt vc_p a_n413_n70# a_n369_101# w_n551_n289# a_n273_n167# VSUBS
X0 a_n273_n167# a_n273_n167# a_n413_n70# w_n551_n289# sky130_fd_pr__pfet_01v8 ad=6.93e+11p pd=6.18e+06u as=1.358e+12p ps=1.228e+07u w=700000u l=150000u
*X1 a_n413_n70# a_n369_101# a_n413_n70# w_n551_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X2 a_n273_n167# a_n273_n167# a_n413_n70# w_n551_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X3 a_n413_n70# a_n273_n167# a_n273_n167# w_n551_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
*X4 a_n413_n70# a_n369_101# a_n413_n70# w_n551_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X5 a_n273_n167# a_n273_n167# a_n413_n70# w_n551_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X6 a_n413_n70# a_n273_n167# a_n273_n167# w_n551_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X7 a_n413_n70# a_n273_n167# a_n273_n167# w_n551_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
C0 a_n413_n70# a_n273_n167# 2.04fF
.ends

.subckt vc_n a_n221_n70# a_n81_92# a_n177_n158# a_n323_n244#
X0 a_n221_n70# a_n81_92# a_n81_92# a_n323_n244# sky130_fd_pr__nfet_01v8 ad=8.96e+11p pd=8.16e+06u as=2.31e+11p ps=2.06e+06u w=700000u l=150000u
X1 a_n81_92# a_n81_92# a_n221_n70# a_n323_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
*X2 a_n221_n70# a_n177_n158# a_n221_n70# a_n323_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
*X3 a_n221_n70# a_n177_n158# a_n221_n70# a_n323_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
.ends

.subckt vc_1 m1_475_n185# sky130_fd_pr__nfet_01v8_2AA63J_0/a_n221_n70# vc_p_0/a_n413_n70#
+ sky130_fd_pr__nfet_01v8_2AA63J_0/a_n177_n158# vc_p_0/a_n369_101# VSUBS vc_p_0/w_n551_n289#
Xvc_p_0 vc_p_0/a_n413_n70# vc_p_0/a_n369_101# vc_p_0/w_n551_n289# m1_475_n185# VSUBS
+ vc_p
Xsky130_fd_pr__nfet_01v8_2AA63J_0 sky130_fd_pr__nfet_01v8_2AA63J_0/a_n221_n70# m1_475_n185#
+ sky130_fd_pr__nfet_01v8_2AA63J_0/a_n177_n158# VSUBS vc_n
C0 vc_p_0/w_n551_n289# VSUBS 2.21fF
.ends

.subckt sinv_p w_n455_n289# a_n317_n70# a_n129_n70# a_n177_n167# a_n273_101# VSUBS
X0 a_n317_n70# a_n177_n167# a_n129_n70# w_n455_n289# sky130_fd_pr__pfet_01v8 ad=1.127e+12p pd=1.022e+07u as=4.62e+11p ps=4.12e+06u w=700000u l=150000u
X1 a_n317_n70# a_n177_n167# a_n129_n70# w_n455_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
*X2 a_n317_n70# a_n273_101# a_n317_n70# w_n455_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
*X3 a_n317_n70# a_n273_101# a_n317_n70# w_n455_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X4 a_n129_n70# a_n177_n167# a_n317_n70# w_n455_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X5 a_n129_n70# a_n177_n167# a_n317_n70# w_n455_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
.ends

.subckt sinv_n a_n221_n70# a_n81_92# a_n33_n70# a_n177_n158# a_n323_n244#
X0 a_n221_n70# a_n81_92# a_n33_n70# a_n323_n244# sky130_fd_pr__nfet_01v8 ad=8.96e+11p pd=8.16e+06u as=2.31e+11p ps=2.06e+06u w=700000u l=150000u
X1 a_n33_n70# a_n81_92# a_n221_n70# a_n323_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
*X2 a_n221_n70# a_n177_n158# a_n221_n70# a_n323_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
*X3 a_n221_n70# a_n177_n158# a_n221_n70# a_n323_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
.ends

.subckt simple_inv m2_381_n263# sky130_fd_pr__nfet_01v8_2AA63J_0/a_n221_n70# sky130_fd_pr__pfet_01v8_X6FFBL_0/w_n455_n289#
+ m1_n53_n74# sky130_fd_pr__nfet_01v8_2AA63J_0/a_n177_n158# sky130_fd_pr__pfet_01v8_X6FFBL_0/a_n317_n70#
+ sky130_fd_pr__pfet_01v8_X6FFBL_0/a_n273_101# VSUBS
Xsky130_fd_pr__pfet_01v8_X6FFBL_0 sky130_fd_pr__pfet_01v8_X6FFBL_0/w_n455_n289# sky130_fd_pr__pfet_01v8_X6FFBL_0/a_n317_n70#
+ m2_381_n263# m1_n53_n74# sky130_fd_pr__pfet_01v8_X6FFBL_0/a_n273_101# VSUBS sinv_p
Xsky130_fd_pr__nfet_01v8_2AA63J_0 sky130_fd_pr__nfet_01v8_2AA63J_0/a_n221_n70# m1_n53_n74#
+ m2_381_n263# sky130_fd_pr__nfet_01v8_2AA63J_0/a_n177_n158# VSUBS sinv_n
.ends

.subckt tg_p a_n221_n70# a_n33_n70# w_n359_n289# a_n81_101# a_n177_n167# VSUBS
X0 a_n33_n70# a_n81_101# a_n221_n70# w_n359_n289# sky130_fd_pr__pfet_01v8 ad=2.31e+11p pd=2.06e+06u as=8.96e+11p ps=8.16e+06u w=700000u l=150000u
*X1 a_n221_n70# a_n177_n167# a_n221_n70# w_n359_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
*X2 a_n221_n70# a_n177_n167# a_n221_n70# w_n359_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X3 a_n221_n70# a_n81_101# a_n33_n70# w_n359_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
.ends

.subckt tg_n a_n221_n70# a_n33_n70# a_n177_92# a_n323_n244# a_n81_n158#
X0 a_n221_n70# a_n81_n158# a_n33_n70# a_n323_n244# sky130_fd_pr__nfet_01v8 ad=8.96e+11p pd=8.16e+06u as=2.31e+11p ps=2.06e+06u w=700000u l=150000u
X1 a_n33_n70# a_n81_n158# a_n221_n70# a_n323_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
*X2 a_n221_n70# a_n177_92# a_n221_n70# a_n323_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
*X3 a_n221_n70# a_n177_92# a_n221_n70# a_n323_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
.ends

.subckt tg_1 sky130_fd_pr__pfet_01v8_X679XQ_0/w_n359_n289# sky130_fd_pr__pfet_01v8_X679XQ_0/a_n81_101#
+ sky130_fd_pr__nfet_01v8_2AA63J_0/a_n177_92# sky130_fd_pr__pfet_01v8_X679XQ_0/a_n177_n167#
+ sky130_fd_pr__nfet_01v8_2AA63J_0/a_n81_n158# m2_477_n333# m2_n53_n74# VSUBS
Xsky130_fd_pr__pfet_01v8_X679XQ_0 m2_477_n333# m2_n53_n74# sky130_fd_pr__pfet_01v8_X679XQ_0/w_n359_n289#
+ sky130_fd_pr__pfet_01v8_X679XQ_0/a_n81_101# sky130_fd_pr__pfet_01v8_X679XQ_0/a_n177_n167#
+ VSUBS tg_p
Xsky130_fd_pr__nfet_01v8_2AA63J_0 m2_477_n333# m2_n53_n74# sky130_fd_pr__nfet_01v8_2AA63J_0/a_n177_92#
+ VSUBS sky130_fd_pr__nfet_01v8_2AA63J_0/a_n81_n158# tg_n
.ends

.subckt tgate_1 m2_717_539# m2_n261_539# simple_inv_0/sky130_fd_pr__pfet_01v8_X6FFBL_0/w_n455_n289#
+ m2_667_n718# m2_0_n814# m1_n261_n952# tg_1_0/sky130_fd_pr__pfet_01v8_X679XQ_0/w_n359_n289#
+ VSUBS
Xsimple_inv_0 m1_282_122# m2_667_n718# simple_inv_0/sky130_fd_pr__pfet_01v8_X6FFBL_0/w_n455_n289#
+ m1_n261_n952# m2_0_n814# m2_0_n814# m2_667_n718# VSUBS simple_inv
Xtg_1_0 tg_1_0/sky130_fd_pr__pfet_01v8_X679XQ_0/w_n359_n289# m1_n261_n952# m2_0_n814#
+ m2_667_n718# m1_282_122# m2_717_539# m2_n261_539# VSUBS tg_1
.ends

.subckt stf_ctrl vdd vss b2 b1 b0 ss tt ff VSUBS
Xvc_1_0 vss vss vdd vdd vss VSUBS vc_1_0/vc_p_0/w_n551_n289# vc_1
Xtgate_1_0 b2 ff tgate_1_1/tg_1_0/sky130_fd_pr__pfet_01v8_X679XQ_0/w_n359_n289# vss
+ vdd vss tgate_1_0/tg_1_0/sky130_fd_pr__pfet_01v8_X679XQ_0/w_n359_n289# VSUBS tgate_1
Xtgate_1_1 b1 tt tgate_1_2/tg_1_0/sky130_fd_pr__pfet_01v8_X679XQ_0/w_n359_n289# vss
+ vdd vss tgate_1_1/tg_1_0/sky130_fd_pr__pfet_01v8_X679XQ_0/w_n359_n289# VSUBS tgate_1
Xtgate_1_2 b0 ss vc_1_0/vc_p_0/w_n551_n289# vss vdd vss tgate_1_2/tg_1_0/sky130_fd_pr__pfet_01v8_X679XQ_0/w_n359_n289#
+ VSUBS tgate_1
C0 vdd VSUBS 6.14fF
C1 vss VSUBS 9.49fF
C2 vc_1_0/vc_p_0/w_n551_n289# VSUBS 3.93fF
C3 tgate_1_2/tg_1_0/sky130_fd_pr__pfet_01v8_X679XQ_0/w_n359_n289# VSUBS 2.88fF
C4 tgate_1_1/tg_1_0/sky130_fd_pr__pfet_01v8_X679XQ_0/w_n359_n289# VSUBS 2.88fF
.ends

.subckt current_tails_2 a_n707_n244# a_n465_n158# a_n561_92# a_n417_n70# a_399_n158#
+ a_n609_n70# a_111_92#
X0 a_n609_n70# a_n465_n158# a_n417_n70# a_n707_n244# sky130_fd_pr__nfet_01v8 ad=1.848e+12p pd=1.648e+07u as=1.155e+12p ps=1.03e+07u w=700000u l=150000u
X1 a_n417_n70# a_n465_n158# a_n609_n70# a_n707_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X2 a_n417_n70# a_111_92# a_n609_n70# a_n707_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X3 a_n609_n70# a_111_92# a_n417_n70# a_n707_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X4 a_n417_n70# a_111_92# a_n609_n70# a_n707_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X5 a_n609_n70# a_399_n158# a_n417_n70# a_n707_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
*X6 a_n609_n70# a_n561_92# a_n609_n70# a_n707_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X7 a_n609_n70# a_n465_n158# a_n417_n70# a_n707_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
*X8 a_n609_n70# a_n561_92# a_n609_n70# a_n707_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X9 a_n417_n70# a_n465_n158# a_n609_n70# a_n707_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X10 a_n417_n70# a_n465_n158# a_n609_n70# a_n707_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X11 a_n609_n70# a_n465_n158# a_n417_n70# a_n707_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
C0 a_n609_n70# a_n417_n70# 4.73fF
.ends

.subckt n_cell a_n321_n70# a_33_n142# a_n419_n244# a_n177_n158# a_63_n70# a_n274_96#
+ a_n129_n70#
X0 a_63_n70# a_33_n142# a_n321_n70# a_n419_n244# sky130_fd_pr__nfet_01v8 ad=2.31e+11p pd=2.06e+06u as=1.155e+12p ps=1.03e+07u w=700000u l=150000u
X1 a_n321_n70# a_n177_n158# a_n129_n70# a_n419_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.31e+11p ps=2.06e+06u w=700000u l=150000u
X2 a_n321_n70# a_33_n142# a_63_n70# a_n419_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
*X3 a_n321_n70# a_n274_96# a_n321_n70# a_n419_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
*X4 a_n321_n70# a_n274_96# a_n321_n70# a_n419_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X5 a_n129_n70# a_n177_n158# a_n321_n70# a_n419_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
.ends

.subckt p_cell_3 a_n321_n70# a_207_n167# a_n369_n167# a_n417_n70# a_303_101# a_n81_101#
+ w_n551_n289# a_n273_101# VSUBS
X0 a_n417_n70# a_n81_101# a_n321_n70# w_n551_n289# sky130_fd_pr__pfet_01v8 ad=1.155e+12p pd=1.03e+07u as=4.62e+11p ps=4.12e+06u w=700000u l=150000u
*X1 a_n417_n70# a_303_101# a_n81_101# w_n551_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.62e+11p ps=4.12e+06u w=700000u l=150000u
X2 a_n417_n70# a_n81_101# a_n81_101# w_n551_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X3 a_n81_101# a_207_n167# a_n417_n70# w_n551_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
*X4 a_n321_n70# a_n369_n167# a_n417_n70# w_n551_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X5 a_n417_n70# a_n273_101# a_n321_n70# w_n551_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X6 a_n321_n70# a_n321_n70# a_n417_n70# w_n551_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X7 a_n81_101# a_n321_n70# a_n417_n70# w_n551_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
.ends

.subckt n_cell_3 a_n32_92# a_n128_n158# a_16_n70# a_n274_n244# a_n172_n70#
X0 a_16_n70# a_n32_92# a_n172_n70# a_n274_n244# sky130_fd_pr__nfet_01v8 ad=2.31e+11p pd=2.06e+06u as=6.79e+11p ps=6.14e+06u w=700000u l=150000u
*X1 a_n172_n70# a_n128_n158# a_n172_n70# a_n274_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
*X2 a_n172_n70# a_n128_n158# a_16_n70# a_n274_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_X679XQ a_n32_n70# a_n80_101# w_n358_n288# a_n176_n167#
+ a_n220_n70# VSUBS
X0 a_n220_n70# a_n80_101# a_n32_n70# w_n358_n288# sky130_fd_pr__pfet_01v8 ad=8.96e+11p pd=8.16e+06u as=2.31e+11p ps=2.06e+06u w=700000u l=150000u
X1 a_n32_n70# a_n80_101# a_n220_n70# w_n358_n288# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
*X2 a_n220_n70# a_n176_n167# a_n220_n70# w_n358_n288# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
*X3 a_n220_n70# a_n176_n167# a_n220_n70# w_n358_n288# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
.ends

.subckt delay_cell_4 sky130_fd_pr__pfet_01v8_X6PFBL_0/w_n551_n289# m2_380_n175# m1_481_490#
+ m1_767_913# m1_863_n597# m1_610_n325# m1_n182_n163# m1_n537_437# m1_707_85# m1_433_n699#
+ m1_n87_n87# m1_920_n163# m2_n115_1015# m3_815_805# VSUBS
Xcurrent_tails_2_0 VSUBS m1_433_n699# m3_815_805# m2_380_n175# m1_863_n597# m1_767_913#
+ m1_610_n325# current_tails_2
Xn_cell_0 m2_380_n175# m1_707_85# VSUBS m1_n87_n87# m1_481_490# m3_815_805# m1_n537_437#
+ n_cell
Xsky130_fd_pr__pfet_01v8_X6PFBL_0 m1_n537_437# m2_n115_1015# m1_767_913# m3_815_805#
+ m1_767_913# m1_481_490# sky130_fd_pr__pfet_01v8_X6PFBL_0/w_n551_n289# m2_n115_1015#
+ VSUBS p_cell_3
Xsky130_fd_pr__nfet_01v8_5ZA63U_0 m1_n537_437# m3_815_805# m1_n182_n163# VSUBS m1_767_913#
+ n_cell_3
Xsky130_fd_pr__nfet_01v8_5ZA63U_1 m1_481_490# m3_815_805# m1_920_n163# VSUBS m1_767_913#
+ n_cell_3
Xsky130_fd_pr__pfet_01v8_X679XQ_0 m1_n182_n163# m1_n537_437# sky130_fd_pr__pfet_01v8_X6PFBL_0/w_n551_n289#
+ m1_767_913# m3_815_805# VSUBS sky130_fd_pr__pfet_01v8_X679XQ
Xsky130_fd_pr__pfet_01v8_X679XQ_1 m1_920_n163# m1_481_490# sky130_fd_pr__pfet_01v8_X6PFBL_0/w_n551_n289#
+ m1_767_913# m3_815_805# VSUBS sky130_fd_pr__pfet_01v8_X679XQ
C0 m3_815_805# VSUBS 3.80fF
C1 m1_767_913# VSUBS 4.07fF
C2 sky130_fd_pr__pfet_01v8_X6PFBL_0/w_n551_n289# VSUBS 5.27fF
.ends

.subckt vco_core_8 inv2 inv1 vdd vss b2 b1 b0 vb2 vb1 out8 out7 out6 out5 out4 out3
+ out2 out1 VSUBS
Xdelay_cell_4_0 delay_cell_4_1/sky130_fd_pr__pfet_01v8_X6PFBL_0/w_n551_n289# m2_1245_n37#
+ out2 vss b2 b1 inv1 out1 out8 b0 out7 inv2 vb2 vdd VSUBS delay_cell_4
Xdelay_cell_4_1 delay_cell_4_1/sky130_fd_pr__pfet_01v8_X6PFBL_0/w_n551_n289# delay_cell_4_1/m2_380_n175#
+ out3 vss b2 b1 inv4 out4 out1 b0 out2 inv3 vb1 vdd VSUBS delay_cell_4
Xdelay_cell_4_2 delay_cell_4_3/sky130_fd_pr__pfet_01v8_X6PFBL_0/w_n551_n289# delay_cell_4_2/m2_380_n175#
+ out6 vss b2 b1 inv5 out5 out3 b0 out4 inv6 vb2 vdd VSUBS delay_cell_4
Xdelay_cell_4_3 delay_cell_4_3/sky130_fd_pr__pfet_01v8_X6PFBL_0/w_n551_n289# delay_cell_4_3/m2_380_n175#
+ out7 vss b2 b1 inv8 out8 out5 b0 out6 inv7 vb1 vdd VSUBS delay_cell_4
*C0 m1_n800_n4112# m1_n1170_n4482# 6.73fF
*C1 m1_n800_n4112# VSUBS 13.30fF **FLOATING
*C2 m1_n1170_n4482# VSUBS 14.90fF **FLOATING
C3 out8 VSUBS 3.78fF
C4 out7 VSUBS 4.46fF
C5 vb1 VSUBS 2.02fF
C6 b2 VSUBS 2.77fF
C7 b0 VSUBS 7.19fF
C8 b1 VSUBS 4.42fF
C9 vss VSUBS 14.56fF
C10 delay_cell_4_3/sky130_fd_pr__pfet_01v8_X6PFBL_0/w_n551_n289# VSUBS 8.77fF
C11 out5 VSUBS 3.92fF
C12 out6 VSUBS 4.32fF
C13 out4 VSUBS 3.49fF
C14 out3 VSUBS 4.53fF
C15 vdd VSUBS 14.06fF
C16 delay_cell_4_1/sky130_fd_pr__pfet_01v8_X6PFBL_0/w_n551_n289# VSUBS 8.77fF
C17 out1 VSUBS 3.49fF
C18 out2 VSUBS 4.60fF
.ends

**.subckt core_complete_1
Xstf_ctrl_0 vdd vss b2 b1 b0 stf_ctrl_0/ss stf_ctrl_0/tt stf_ctrl_0/ff VSUBS stf_ctrl
Xvco_core_8_0 inv2 inv1 vdd vss b2 b1 b0 vb2 vb1 vco_core_8_0/out8 vco_core_8_0/out7
+ vco_core_8_0/out6 vco_core_8_0/out5 vco_core_8_0/out4 vco_core_8_0/out3 out2 out1
+ VSUBS vco_core_8
C0 b1 b2 9.04fF
C1 b1 b0 6.84fF
C2 b0 b2 2.70fF
*C3 vco_core_8_0/m1_n800_n4112# VSUBS 13.30fF **FLOATING
*C4 vco_core_8_0/m1_n1170_n4482# VSUBS 14.90fF **FLOATING
C5 vco_core_8_0/out8 VSUBS 3.72fF
C6 vco_core_8_0/out7 VSUBS 4.40fF
C7 vb1 VSUBS 2.32fF
C8 b2 VSUBS 6.37fF
C9 b0 VSUBS 9.63fF
C10 b1 VSUBS 7.15fF
C11 vss VSUBS 24.40fF
*C12 vco_core_8_0/delay_cell_4_3/sky130_fd_pr__pfet_01v8_X6PFBL_0/w_n551_n289# VSUBS 8.77fF
C13 vco_core_8_0/out5 VSUBS 3.86fF
C14 vco_core_8_0/out6 VSUBS 4.32fF
C15 vco_core_8_0/out4 VSUBS 3.25fF
C16 vco_core_8_0/out3 VSUBS 4.37fF
C17 vdd VSUBS 20.51fF
*C18 vco_core_8_0/delay_cell_4_1/sky130_fd_pr__pfet_01v8_X6PFBL_0/w_n551_n289# VSUBS 8.77fF
C19 out1 VSUBS 3.69fF
C20 out2 VSUBS 4.75fF
*C21 stf_ctrl_0/vc_1_0/vc_p_0/w_n551_n289# VSUBS 3.93fF
*C22 stf_ctrl_0/tgate_1_2/tg_1_0/sky130_fd_pr__pfet_01v8_X679XQ_0/w_n359_n289# VSUBS 2.82fF
*C23 stf_ctrl_0/tgate_1_1/tg_1_0/sky130_fd_pr__pfet_01v8_X679XQ_0/w_n359_n289# VSUBS 2.82fF
**.ends
**** begin user architecture code

.lib /foss/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice.tt.red tt

.control
set temp=25
alter v10 1.8
alter v11 0
alter v12 1.8
save out1 out2 inv1 inv2 @V4[i]
tran 0.01n 100n 50n
plot out1 out2
fft out1 inv1
plot db(mag(out1)) db(mag(inv1)) xlimit 0.5g 10g ylimit 0.0 -200
.endc
.end

**** end user architecture code
