magic
tech sky130A
magscale 1 2
timestamp 1663426905
<< error_p >>
rect -557 151 -499 157
rect 499 151 557 157
rect -557 117 -545 151
rect 499 117 511 151
rect -557 111 -499 117
rect 499 111 557 117
<< nwell >>
rect -743 -289 743 289
<< pmos >>
rect -543 -70 -513 70
rect -447 -70 -417 70
rect -351 -70 -321 70
rect -255 -70 -225 70
rect -159 -70 -129 70
rect -63 -70 -33 70
rect 33 -70 63 70
rect 129 -70 159 70
rect 225 -70 255 70
rect 321 -70 351 70
rect 417 -70 447 70
rect 513 -70 543 70
<< pdiff >>
rect -605 58 -543 70
rect -605 -58 -593 58
rect -559 -58 -543 58
rect -605 -70 -543 -58
rect -513 58 -447 70
rect -513 -58 -497 58
rect -463 -58 -447 58
rect -513 -70 -447 -58
rect -417 58 -351 70
rect -417 -58 -401 58
rect -367 -58 -351 58
rect -417 -70 -351 -58
rect -321 58 -255 70
rect -321 -58 -305 58
rect -271 -58 -255 58
rect -321 -70 -255 -58
rect -225 58 -159 70
rect -225 -58 -209 58
rect -175 -58 -159 58
rect -225 -70 -159 -58
rect -129 58 -63 70
rect -129 -58 -113 58
rect -79 -58 -63 58
rect -129 -70 -63 -58
rect -33 58 33 70
rect -33 -58 -17 58
rect 17 -58 33 58
rect -33 -70 33 -58
rect 63 58 129 70
rect 63 -58 79 58
rect 113 -58 129 58
rect 63 -70 129 -58
rect 159 58 225 70
rect 159 -58 175 58
rect 209 -58 225 58
rect 159 -70 225 -58
rect 255 58 321 70
rect 255 -58 271 58
rect 305 -58 321 58
rect 255 -70 321 -58
rect 351 58 417 70
rect 351 -58 367 58
rect 401 -58 417 58
rect 351 -70 417 -58
rect 447 58 513 70
rect 447 -58 463 58
rect 497 -58 513 58
rect 447 -70 513 -58
rect 543 58 609 70
rect 543 -58 559 58
rect 593 -2 609 58
rect 593 -58 605 -2
rect 543 -70 605 -58
<< pdiffc >>
rect -593 -58 -559 58
rect -497 -58 -463 58
rect -401 -58 -367 58
rect -305 -58 -271 58
rect -209 -58 -175 58
rect -113 -58 -79 58
rect -17 -58 17 58
rect 79 -58 113 58
rect 175 -58 209 58
rect 271 -58 305 58
rect 367 -58 401 58
rect 463 -58 497 58
rect 559 -58 593 58
<< nsubdiff >>
rect -707 219 -611 253
rect 611 219 707 253
rect -707 157 -673 219
rect 673 157 707 219
rect -707 -219 -673 -157
rect 673 -219 707 -157
rect -707 -253 -611 -219
rect 611 -253 707 -219
<< nsubdiffcont >>
rect -611 219 611 253
rect -707 -157 -673 157
rect 673 -157 707 157
rect -611 -253 611 -219
<< poly >>
rect -561 151 -495 167
rect -561 117 -545 151
rect -511 117 -495 151
rect -561 101 -495 117
rect 495 151 561 167
rect 495 117 511 151
rect 545 117 561 151
rect 495 101 561 117
rect -543 70 -513 101
rect -447 70 -417 96
rect -351 70 -321 96
rect -255 70 -225 96
rect -159 70 -129 96
rect -63 70 -33 96
rect 33 70 63 96
rect 129 70 159 96
rect 225 70 255 96
rect 321 70 351 96
rect 417 70 447 96
rect 513 70 543 101
rect -543 -96 -513 -70
rect -447 -101 -417 -70
rect -351 -101 -321 -70
rect -255 -101 -225 -70
rect -159 -101 -129 -70
rect -63 -101 -33 -70
rect 33 -101 63 -70
rect 129 -101 159 -70
rect 225 -101 255 -70
rect 321 -101 351 -70
rect 417 -101 447 -70
rect 513 -96 543 -70
rect -465 -117 465 -101
rect -465 -151 -449 -117
rect -415 -151 -353 -117
rect -319 -151 -257 -117
rect -223 -151 -161 -117
rect -127 -151 -65 -117
rect -31 -151 31 -117
rect 65 -151 127 -117
rect 161 -151 223 -117
rect 257 -151 319 -117
rect 353 -151 415 -117
rect 449 -151 465 -117
rect -465 -167 465 -151
<< polycont >>
rect -545 117 -511 151
rect 511 117 545 151
rect -449 -151 -415 -117
rect -353 -151 -319 -117
rect -257 -151 -223 -117
rect -161 -151 -127 -117
rect -65 -151 -31 -117
rect 31 -151 65 -117
rect 127 -151 161 -117
rect 223 -151 257 -117
rect 319 -151 353 -117
rect 415 -151 449 -117
<< locali >>
rect -707 219 -611 253
rect 611 219 707 253
rect -707 157 -673 219
rect 673 157 707 219
rect -561 117 -545 151
rect -511 117 -495 151
rect 495 117 511 151
rect 545 117 561 151
rect -593 58 -559 74
rect -593 -74 -559 -58
rect -497 58 -463 74
rect -497 -74 -463 -58
rect -401 58 -367 74
rect -401 -74 -367 -58
rect -305 58 -271 74
rect -305 -74 -271 -58
rect -209 58 -175 74
rect -209 -74 -175 -58
rect -113 58 -79 74
rect -113 -74 -79 -58
rect -17 58 17 74
rect -17 -74 17 -58
rect 79 58 113 74
rect 79 -74 113 -58
rect 175 58 209 74
rect 175 -74 209 -58
rect 271 58 305 74
rect 271 -74 305 -58
rect 367 58 401 74
rect 367 -74 401 -58
rect 463 58 497 74
rect 463 -74 497 -58
rect 559 58 593 74
rect 559 -74 593 -58
rect -465 -151 -449 -117
rect -415 -151 -353 -117
rect -319 -151 -257 -117
rect -223 -151 -161 -117
rect -127 -151 -65 -117
rect -31 -151 31 -117
rect 65 -151 127 -117
rect 161 -151 223 -117
rect 257 -151 319 -117
rect 353 -151 415 -117
rect 449 -151 465 -117
rect -707 -219 -673 -157
rect 673 -219 707 -157
rect -707 -253 -611 -219
rect 611 -253 707 -219
<< viali >>
rect -545 117 -511 151
rect 511 117 545 151
rect -593 -58 -559 58
rect -497 -58 -463 58
rect -401 -58 -367 58
rect -305 -58 -271 58
rect -209 -58 -175 58
rect -113 -58 -79 58
rect -17 -58 17 58
rect 79 -58 113 58
rect 175 -58 209 58
rect 271 -58 305 58
rect 367 -58 401 58
rect 463 -58 497 58
rect 559 -58 593 58
rect -449 -151 -415 -117
rect -353 -151 -319 -117
rect -257 -151 -223 -117
rect -161 -151 -127 -117
rect -65 -151 -31 -117
rect 31 -151 65 -117
rect 127 -151 161 -117
rect 223 -151 257 -117
rect 319 -151 353 -117
rect 415 -151 449 -117
<< metal1 >>
rect -557 151 -499 157
rect -557 117 -545 151
rect -511 117 -499 151
rect -557 111 -499 117
rect 499 151 557 157
rect 499 117 511 151
rect 545 117 557 151
rect 499 111 557 117
rect -607 61 -545 70
rect -607 9 -602 61
rect -550 9 -545 61
rect -607 0 -593 9
rect -599 -58 -593 0
rect -559 0 -545 9
rect -511 61 -449 70
rect -511 9 -506 61
rect -454 9 -449 61
rect -511 0 -497 9
rect -559 -58 -553 0
rect -599 -70 -553 -58
rect -503 -58 -497 0
rect -463 0 -449 9
rect -407 58 -361 70
rect -407 0 -401 58
rect -463 -58 -457 0
rect -503 -70 -457 -58
rect -415 -9 -401 0
rect -367 0 -361 58
rect -319 61 -257 70
rect -319 9 -314 61
rect -262 9 -257 61
rect -319 0 -305 9
rect -367 -9 -353 0
rect -415 -61 -410 -9
rect -358 -61 -353 -9
rect -415 -70 -353 -61
rect -311 -58 -305 0
rect -271 0 -257 9
rect -215 58 -169 70
rect -215 0 -209 58
rect -271 -58 -265 0
rect -311 -70 -265 -58
rect -223 -9 -209 0
rect -175 0 -169 58
rect -127 61 -65 70
rect -127 9 -122 61
rect -70 9 -65 61
rect -127 0 -113 9
rect -175 -9 -161 0
rect -223 -61 -218 -9
rect -166 -61 -161 -9
rect -223 -70 -161 -61
rect -119 -58 -113 0
rect -79 0 -65 9
rect -23 58 23 70
rect -23 0 -17 58
rect -79 -58 -73 0
rect -119 -70 -73 -58
rect -31 -9 -17 0
rect 17 0 23 58
rect 65 61 127 70
rect 65 9 70 61
rect 122 9 127 61
rect 65 0 79 9
rect 17 -9 31 0
rect -31 -61 -26 -9
rect 26 -61 31 -9
rect -31 -70 31 -61
rect 73 -58 79 0
rect 113 0 127 9
rect 169 58 215 70
rect 169 0 175 58
rect 113 -58 119 0
rect 73 -70 119 -58
rect 161 -9 175 0
rect 209 0 215 58
rect 257 61 319 70
rect 257 9 262 61
rect 314 9 319 61
rect 257 0 271 9
rect 209 -9 223 0
rect 161 -61 166 -9
rect 218 -61 223 -9
rect 161 -70 223 -61
rect 265 -58 271 0
rect 305 0 319 9
rect 361 58 407 70
rect 361 0 367 58
rect 305 -58 311 0
rect 265 -70 311 -58
rect 353 -9 367 0
rect 401 0 407 58
rect 449 61 511 70
rect 449 9 454 61
rect 506 9 511 61
rect 449 0 463 9
rect 401 -9 415 0
rect 353 -61 358 -9
rect 410 -61 415 -9
rect 353 -70 415 -61
rect 457 -58 463 0
rect 497 0 511 9
rect 545 61 607 70
rect 545 9 550 61
rect 602 9 607 61
rect 545 0 559 9
rect 497 -58 503 0
rect 457 -70 503 -58
rect 553 -58 559 0
rect 593 0 607 9
rect 593 -58 599 0
rect 553 -70 599 -58
rect -461 -117 -403 -111
rect -365 -117 -307 -111
rect -269 -117 -211 -111
rect -173 -117 -115 -111
rect -77 -117 -19 -111
rect 19 -117 77 -111
rect 115 -117 173 -111
rect 211 -117 269 -111
rect 307 -117 365 -111
rect 403 -117 461 -111
rect -461 -151 -449 -117
rect -415 -151 -353 -117
rect -319 -151 -257 -117
rect -223 -151 -161 -117
rect -127 -151 -65 -117
rect -31 -151 31 -117
rect 65 -151 127 -117
rect 161 -151 223 -117
rect 257 -151 319 -117
rect 353 -151 415 -117
rect 449 -151 461 -117
rect -461 -157 -403 -151
rect -365 -157 -307 -151
rect -269 -157 -211 -151
rect -173 -157 -115 -151
rect -77 -157 -19 -151
rect 19 -157 77 -151
rect 115 -157 173 -151
rect 211 -157 269 -151
rect 307 -157 365 -151
rect 403 -157 461 -151
<< via1 >>
rect -602 58 -550 61
rect -602 9 -593 58
rect -593 9 -559 58
rect -559 9 -550 58
rect -506 58 -454 61
rect -506 9 -497 58
rect -497 9 -463 58
rect -463 9 -454 58
rect -314 58 -262 61
rect -314 9 -305 58
rect -305 9 -271 58
rect -271 9 -262 58
rect -410 -58 -401 -9
rect -401 -58 -367 -9
rect -367 -58 -358 -9
rect -410 -61 -358 -58
rect -122 58 -70 61
rect -122 9 -113 58
rect -113 9 -79 58
rect -79 9 -70 58
rect -218 -58 -209 -9
rect -209 -58 -175 -9
rect -175 -58 -166 -9
rect -218 -61 -166 -58
rect 70 58 122 61
rect 70 9 79 58
rect 79 9 113 58
rect 113 9 122 58
rect -26 -58 -17 -9
rect -17 -58 17 -9
rect 17 -58 26 -9
rect -26 -61 26 -58
rect 262 58 314 61
rect 262 9 271 58
rect 271 9 305 58
rect 305 9 314 58
rect 166 -58 175 -9
rect 175 -58 209 -9
rect 209 -58 218 -9
rect 166 -61 218 -58
rect 454 58 506 61
rect 454 9 463 58
rect 463 9 497 58
rect 497 9 506 58
rect 358 -58 367 -9
rect 367 -58 401 -9
rect 401 -58 410 -9
rect 358 -61 410 -58
rect 550 58 602 61
rect 550 9 559 58
rect 559 9 593 58
rect 593 9 602 58
<< metal2 >>
rect -613 63 -443 72
rect -613 7 -604 63
rect -548 7 -508 63
rect -452 7 -443 63
rect -613 -2 -443 7
rect -325 63 -251 72
rect -325 7 -316 63
rect -260 7 -251 63
rect -415 -9 -353 0
rect -325 -2 -251 7
rect -133 63 -59 72
rect -133 7 -124 63
rect -68 7 -59 63
rect -415 -61 -410 -9
rect -358 -36 -353 -9
rect -223 -9 -161 0
rect -133 -2 -59 7
rect 59 63 133 72
rect 59 7 68 63
rect 124 7 133 63
rect -223 -36 -218 -9
rect -358 -61 -218 -36
rect -166 -36 -161 -9
rect -31 -9 31 0
rect 59 -2 133 7
rect 251 63 325 72
rect 251 7 260 63
rect 316 7 325 63
rect -31 -36 -26 -9
rect -166 -61 -26 -36
rect 26 -36 31 -9
rect 161 -9 223 0
rect 251 -2 325 7
rect 443 63 613 72
rect 443 7 452 63
rect 508 7 548 63
rect 604 7 613 63
rect 161 -36 166 -9
rect 26 -61 166 -36
rect 218 -36 223 -9
rect 353 -9 415 0
rect 443 -2 613 7
rect 353 -36 358 -9
rect 218 -61 358 -36
rect 410 -61 415 -9
rect -415 -70 415 -61
<< via2 >>
rect -604 61 -548 63
rect -604 9 -602 61
rect -602 9 -550 61
rect -550 9 -548 61
rect -604 7 -548 9
rect -508 61 -452 63
rect -508 9 -506 61
rect -506 9 -454 61
rect -454 9 -452 61
rect -508 7 -452 9
rect -316 61 -260 63
rect -316 9 -314 61
rect -314 9 -262 61
rect -262 9 -260 61
rect -316 7 -260 9
rect -124 61 -68 63
rect -124 9 -122 61
rect -122 9 -70 61
rect -70 9 -68 61
rect -124 7 -68 9
rect 68 61 124 63
rect 68 9 70 61
rect 70 9 122 61
rect 122 9 124 61
rect 68 7 124 9
rect 260 61 316 63
rect 260 9 262 61
rect 262 9 314 61
rect 314 9 316 61
rect 260 7 316 9
rect 452 61 508 63
rect 452 9 454 61
rect 454 9 506 61
rect 506 9 508 61
rect 452 7 508 9
rect 548 61 604 63
rect 548 9 550 61
rect 550 9 602 61
rect 602 9 604 61
rect 548 7 604 9
<< metal3 >>
rect -613 70 -443 72
rect -325 70 -251 72
rect -133 70 -59 72
rect 59 70 133 72
rect 251 70 325 72
rect 443 70 613 72
rect -613 63 613 70
rect -613 7 -604 63
rect -548 7 -508 63
rect -452 10 -316 63
rect -452 7 -443 10
rect -613 -2 -443 7
rect -325 7 -316 10
rect -260 10 -124 63
rect -260 7 -251 10
rect -325 -2 -251 7
rect -133 7 -124 10
rect -68 10 68 63
rect -68 7 -59 10
rect -133 -2 -59 7
rect 59 7 68 10
rect 124 10 260 63
rect 124 7 133 10
rect 59 -2 133 7
rect 251 7 260 10
rect 316 10 452 63
rect 316 7 325 10
rect 251 -2 325 7
rect 443 7 452 10
rect 508 7 548 63
rect 604 7 613 63
rect 443 -2 613 7
<< properties >>
string FIXED_BBOX -690 -236 690 236
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.7 l 0.15 m 1 nf 12 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
