magic
tech sky130A
magscale 1 2
timestamp 1660924145
<< nwell >>
rect -551 -289 551 289
<< pmos >>
rect -351 -70 -321 70
rect -255 -70 -225 70
rect -159 -70 -129 70
rect -63 -70 -33 70
rect 33 -70 63 70
rect 129 -70 159 70
rect 225 -70 255 70
rect 321 -70 351 70
<< pdiff >>
rect -413 58 -351 70
rect -413 -58 -401 58
rect -367 -58 -351 58
rect -413 -70 -351 -58
rect -321 58 -255 70
rect -321 -58 -305 58
rect -271 -58 -255 58
rect -321 -70 -255 -58
rect -225 58 -159 70
rect -225 -58 -209 58
rect -175 -58 -159 58
rect -225 -70 -159 -58
rect -129 58 -63 70
rect -129 -58 -113 58
rect -79 -58 -63 58
rect -129 -70 -63 -58
rect -33 58 33 70
rect -33 -58 -17 58
rect 17 -58 33 58
rect -33 -70 33 -58
rect 63 58 129 70
rect 63 -58 79 58
rect 113 -58 129 58
rect 63 -70 129 -58
rect 159 58 225 70
rect 159 -58 175 58
rect 209 -58 225 58
rect 159 -70 225 -58
rect 255 58 321 70
rect 255 -58 271 58
rect 305 -58 321 58
rect 255 -70 321 -58
rect 351 58 413 70
rect 351 -58 367 58
rect 401 -58 413 58
rect 351 -70 413 -58
<< pdiffc >>
rect -401 -58 -367 58
rect -305 -58 -271 58
rect -209 -58 -175 58
rect -113 -58 -79 58
rect -17 -58 17 58
rect 79 -58 113 58
rect 175 -58 209 58
rect 271 -58 305 58
rect 367 -58 401 58
<< nsubdiff >>
rect -515 219 -419 253
rect 419 219 515 253
rect -515 157 -481 219
rect 481 157 515 219
rect -515 -219 -481 -157
rect 481 -219 515 -157
rect -515 -253 -419 -219
rect 419 -253 515 -219
<< nsubdiffcont >>
rect -419 219 419 253
rect -515 -157 -481 157
rect 481 -157 515 157
rect -419 -253 419 -219
<< poly >>
rect -369 151 -303 167
rect -369 117 -353 151
rect -319 117 -303 151
rect -369 101 -303 117
rect 303 151 369 167
rect 303 117 319 151
rect 353 117 369 151
rect 303 101 369 117
rect -351 70 -321 101
rect -255 70 -225 96
rect -159 70 -129 96
rect -63 70 -33 96
rect 33 70 63 96
rect 129 70 159 96
rect 225 70 255 96
rect 321 70 351 101
rect -351 -96 -321 -70
rect -255 -101 -225 -70
rect -159 -101 -129 -70
rect -63 -101 -33 -70
rect 33 -101 63 -70
rect 129 -101 159 -70
rect 225 -101 255 -70
rect 321 -96 351 -70
rect -273 -117 273 -101
rect -273 -151 -257 -117
rect -223 -151 -161 -117
rect -127 -151 -65 -117
rect -31 -151 31 -117
rect 65 -151 127 -117
rect 161 -151 223 -117
rect 257 -151 273 -117
rect -273 -167 273 -151
<< polycont >>
rect -353 117 -319 151
rect 319 117 353 151
rect -257 -151 -223 -117
rect -161 -151 -127 -117
rect -65 -151 -31 -117
rect 31 -151 65 -117
rect 127 -151 161 -117
rect 223 -151 257 -117
<< locali >>
rect -515 219 -419 253
rect 419 219 515 253
rect -515 157 -481 219
rect 481 157 515 219
rect -369 117 -353 151
rect -319 117 -303 151
rect 303 117 319 151
rect 353 117 369 151
rect -401 58 -367 74
rect -401 -74 -367 -58
rect -305 58 -271 74
rect -305 -74 -271 -58
rect -209 58 -175 74
rect -209 -74 -175 -58
rect -113 58 -79 74
rect -113 -74 -79 -58
rect -17 58 17 74
rect -17 -74 17 -58
rect 79 58 113 74
rect 79 -74 113 -58
rect 175 58 209 74
rect 175 -74 209 -58
rect 271 58 305 74
rect 271 -74 305 -58
rect 367 58 401 74
rect 367 -74 401 -58
rect -273 -151 -257 -117
rect -223 -151 -161 -117
rect -127 -151 -65 -117
rect -31 -151 31 -117
rect 65 -151 127 -117
rect 161 -151 223 -117
rect 257 -151 273 -117
rect -515 -219 -481 -157
rect 481 -219 515 -157
rect -515 -253 -419 -219
rect 419 -253 515 -219
<< viali >>
rect -353 117 -319 151
rect 319 117 353 151
rect -401 -58 -367 58
rect -305 -58 -271 58
rect -209 -58 -175 58
rect -113 -58 -79 58
rect -17 -58 17 58
rect 79 -58 113 58
rect 175 -58 209 58
rect 271 -58 305 58
rect 367 -58 401 58
rect -257 -151 -223 -117
rect -161 -151 -127 -117
rect -65 -151 -31 -117
rect 31 -151 65 -117
rect 127 -151 161 -117
rect 223 -151 257 -117
<< metal1 >>
rect -365 151 -307 157
rect 307 151 365 157
rect -365 117 -353 151
rect -319 117 319 151
rect 353 117 365 151
rect -365 111 -307 117
rect 307 111 365 117
rect -413 60 -259 70
rect -413 8 -410 60
rect -358 8 -314 60
rect -262 8 -259 60
rect -413 0 -401 8
rect -407 -58 -401 0
rect -367 0 -305 8
rect -367 -58 -361 0
rect -407 -70 -361 -58
rect -311 -58 -305 0
rect -271 0 -259 8
rect -215 58 -169 70
rect -271 -58 -265 0
rect -311 -70 -265 -58
rect -215 -58 -209 58
rect -175 -58 -169 58
rect -125 60 -67 70
rect -125 8 -122 60
rect -70 8 -67 60
rect -125 0 -113 8
rect -215 -111 -169 -58
rect -119 -58 -113 0
rect -79 0 -67 8
rect -23 58 23 70
rect -79 -58 -73 0
rect -119 -70 -73 -58
rect -23 -58 -17 58
rect 17 -58 23 58
rect 67 60 125 70
rect 67 8 70 60
rect 122 8 125 60
rect 67 0 79 8
rect -23 -111 23 -58
rect 73 -58 79 0
rect 113 0 125 8
rect 169 58 215 70
rect 113 -58 119 0
rect 73 -70 119 -58
rect 169 -58 175 58
rect 209 -58 215 58
rect 259 60 413 70
rect 259 8 262 60
rect 314 8 358 60
rect 410 8 413 60
rect 259 0 271 8
rect 169 -111 215 -58
rect 265 -58 271 0
rect 305 0 367 8
rect 305 -58 311 0
rect 265 -70 311 -58
rect 361 -58 367 0
rect 401 0 413 8
rect 401 -58 407 0
rect 361 -70 407 -58
rect -269 -117 269 -111
rect -269 -151 -257 -117
rect -223 -151 -161 -117
rect -127 -151 -65 -117
rect -31 -151 31 -117
rect 65 -151 127 -117
rect 161 -151 223 -117
rect 257 -151 269 -117
rect -269 -157 269 -151
<< via1 >>
rect -410 58 -358 60
rect -410 8 -401 58
rect -401 8 -367 58
rect -367 8 -358 58
rect -314 58 -262 60
rect -314 8 -305 58
rect -305 8 -271 58
rect -271 8 -262 58
rect -122 58 -70 60
rect -122 8 -113 58
rect -113 8 -79 58
rect -79 8 -70 58
rect 70 58 122 60
rect 70 8 79 58
rect 79 8 113 58
rect 113 8 122 58
rect 262 58 314 60
rect 262 8 271 58
rect 271 8 305 58
rect 305 8 314 58
rect 358 58 410 60
rect 358 8 367 58
rect 367 8 401 58
rect 401 8 410 58
<< metal2 >>
rect -413 60 413 70
rect -413 8 -410 60
rect -358 8 -314 60
rect -262 28 -122 60
rect -262 8 -259 28
rect -413 0 -259 8
rect -125 8 -122 28
rect -70 28 70 60
rect -70 8 -67 28
rect -125 0 -67 8
rect 67 8 70 28
rect 122 28 262 60
rect 122 8 125 28
rect 67 0 125 8
rect 259 8 262 28
rect 314 8 358 60
rect 410 8 413 60
rect 259 0 413 8
<< properties >>
string FIXED_BBOX -498 -236 498 236
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.7 l 0.15 m 1 nf 8 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
