magic
tech sky130A
magscale 1 2
timestamp 1667124946
<< error_p >>
rect 595 142 653 148
rect 595 108 607 142
rect 595 102 653 108
rect -653 -108 -595 -102
rect -653 -142 -641 -108
rect -653 -148 -595 -142
<< pwell >>
rect -839 -280 839 280
<< nmos >>
rect -639 -70 -609 70
rect -543 -70 -513 70
rect -447 -70 -417 70
rect -351 -70 -321 70
rect -255 -70 -225 70
rect -159 -70 -129 70
rect -63 -70 -33 70
rect 33 -70 63 70
rect 129 -70 159 70
rect 225 -70 255 70
rect 321 -70 351 70
rect 417 -70 447 70
rect 513 -70 543 70
rect 609 -70 639 70
<< ndiff >>
rect -701 58 -639 70
rect -701 -58 -689 58
rect -655 -58 -639 58
rect -701 -70 -639 -58
rect -609 58 -543 70
rect -609 -58 -593 58
rect -559 -58 -543 58
rect -609 -70 -543 -58
rect -513 58 -447 70
rect -513 -58 -497 58
rect -463 -58 -447 58
rect -513 -70 -447 -58
rect -417 58 -351 70
rect -417 -58 -401 58
rect -367 -58 -351 58
rect -417 -70 -351 -58
rect -321 58 -255 70
rect -321 -58 -305 58
rect -271 -58 -255 58
rect -321 -70 -255 -58
rect -225 58 -159 70
rect -225 -58 -209 58
rect -175 -58 -159 58
rect -225 -70 -159 -58
rect -129 58 -63 70
rect -129 -58 -113 58
rect -79 -58 -63 58
rect -129 -70 -63 -58
rect -33 58 33 70
rect -33 -58 -17 58
rect 17 -58 33 58
rect -33 -70 33 -58
rect 63 58 129 70
rect 63 -58 79 58
rect 113 -58 129 58
rect 63 -70 129 -58
rect 159 58 225 70
rect 159 -58 175 58
rect 209 -58 225 58
rect 159 -70 225 -58
rect 255 58 321 70
rect 255 -58 271 58
rect 305 -58 321 58
rect 255 -70 321 -58
rect 351 58 417 70
rect 351 -58 367 58
rect 401 -58 417 58
rect 351 -70 417 -58
rect 447 58 513 70
rect 447 -58 463 58
rect 497 -58 513 58
rect 447 -70 513 -58
rect 543 58 609 70
rect 543 -58 559 58
rect 593 -58 609 58
rect 543 -70 609 -58
rect 639 58 701 70
rect 639 -58 655 58
rect 689 -58 701 58
rect 639 -70 701 -58
<< ndiffc >>
rect -689 -58 -655 58
rect -593 -58 -559 58
rect -497 -58 -463 58
rect -401 -58 -367 58
rect -305 -58 -271 58
rect -209 -58 -175 58
rect -113 -58 -79 58
rect -17 -58 17 58
rect 79 -58 113 58
rect 175 -58 209 58
rect 271 -58 305 58
rect 367 -58 401 58
rect 463 -58 497 58
rect 559 -58 593 58
rect 655 -58 689 58
<< psubdiff >>
rect -803 210 -707 244
rect 707 210 803 244
rect -803 148 -769 210
rect 769 148 803 210
rect -803 -210 -769 -148
rect 769 -210 803 -148
rect -803 -244 -707 -210
rect 707 -244 803 -210
<< psubdiffcont >>
rect -707 210 707 244
rect -803 -148 -769 148
rect 769 -148 803 148
rect -707 -244 707 -210
<< poly >>
rect -561 142 369 158
rect -561 108 -545 142
rect -511 108 -449 142
rect -415 108 -353 142
rect -319 108 -257 142
rect -223 108 -161 142
rect -127 108 -65 142
rect -31 108 31 142
rect 65 108 127 142
rect 161 108 223 142
rect 257 108 319 142
rect 353 108 369 142
rect -639 70 -609 96
rect -561 92 369 108
rect 591 142 657 158
rect 591 108 607 142
rect 641 108 657 142
rect -543 70 -513 92
rect -447 70 -417 92
rect -351 70 -321 92
rect -255 70 -225 92
rect -159 70 -129 92
rect -63 70 -33 92
rect 33 70 63 92
rect 129 70 159 92
rect 225 70 255 92
rect 321 70 351 92
rect 417 70 447 96
rect 513 70 543 96
rect 591 92 657 108
rect 609 70 639 92
rect -639 -92 -609 -70
rect -657 -108 -591 -92
rect -543 -96 -513 -70
rect -447 -96 -417 -70
rect -351 -96 -321 -70
rect -255 -96 -225 -70
rect -159 -96 -129 -70
rect -63 -96 -33 -70
rect 33 -96 63 -70
rect 129 -96 159 -70
rect 225 -96 255 -70
rect 321 -96 351 -70
rect 417 -92 447 -70
rect 513 -92 543 -70
rect -657 -142 -641 -108
rect -607 -142 -591 -108
rect -657 -158 -591 -142
rect 399 -108 561 -92
rect 609 -96 639 -70
rect 399 -142 415 -108
rect 449 -142 511 -108
rect 545 -142 561 -108
rect 399 -158 561 -142
<< polycont >>
rect -545 108 -511 142
rect -449 108 -415 142
rect -353 108 -319 142
rect -257 108 -223 142
rect -161 108 -127 142
rect -65 108 -31 142
rect 31 108 65 142
rect 127 108 161 142
rect 223 108 257 142
rect 319 108 353 142
rect 607 108 641 142
rect -641 -142 -607 -108
rect 415 -142 449 -108
rect 511 -142 545 -108
<< locali >>
rect -803 210 -707 244
rect 707 210 803 244
rect -803 148 -769 210
rect 769 148 803 210
rect -561 108 -545 142
rect -511 108 -449 142
rect -415 108 -353 142
rect -319 108 -257 142
rect -223 108 -161 142
rect -127 108 -65 142
rect -31 108 31 142
rect 65 108 127 142
rect 161 108 223 142
rect 257 108 319 142
rect 353 108 369 142
rect 591 108 607 142
rect 641 108 657 142
rect -689 58 -655 74
rect -689 -74 -655 -58
rect -593 58 -559 74
rect -593 -74 -559 -58
rect -497 58 -463 74
rect -497 -74 -463 -58
rect -401 58 -367 74
rect -401 -74 -367 -58
rect -305 58 -271 74
rect -305 -74 -271 -58
rect -209 58 -175 74
rect -209 -74 -175 -58
rect -113 58 -79 74
rect -113 -74 -79 -58
rect -17 58 17 74
rect -17 -74 17 -58
rect 79 58 113 74
rect 79 -74 113 -58
rect 175 58 209 74
rect 175 -74 209 -58
rect 271 58 305 74
rect 271 -74 305 -58
rect 367 58 401 74
rect 367 -74 401 -58
rect 463 58 497 74
rect 463 -74 497 -58
rect 559 58 593 74
rect 559 -74 593 -58
rect 655 58 689 74
rect 655 -74 689 -58
rect -657 -142 -641 -108
rect -607 -142 -591 -108
rect 399 -142 415 -108
rect 449 -142 511 -108
rect 545 -142 561 -108
rect -803 -210 -769 -148
rect 769 -210 803 -148
rect -803 -244 -707 -210
rect 707 -244 803 -210
<< viali >>
rect -545 108 -511 142
rect -449 108 -415 142
rect -353 108 -319 142
rect -257 108 -223 142
rect -161 108 -127 142
rect -65 108 -31 142
rect 31 108 65 142
rect 127 108 161 142
rect 223 108 257 142
rect 319 108 353 142
rect 607 108 641 142
rect -689 -58 -655 58
rect -593 -58 -559 58
rect -497 -58 -463 58
rect -401 -58 -367 58
rect -305 -58 -271 58
rect -209 -58 -175 58
rect -113 -58 -79 58
rect -17 -58 17 58
rect 79 -58 113 58
rect 175 -58 209 58
rect 271 -58 305 58
rect 367 -58 401 58
rect 463 -58 497 58
rect 559 -58 593 58
rect 655 -58 689 58
rect -641 -142 -607 -108
rect 415 -142 449 -108
rect 511 -142 545 -108
<< metal1 >>
rect -561 142 369 149
rect -561 108 -545 142
rect -511 108 -449 142
rect -415 108 -353 142
rect -319 108 -257 142
rect -223 108 -161 142
rect -127 108 -65 142
rect -31 108 31 142
rect 65 108 127 142
rect 161 108 223 142
rect 257 108 319 142
rect 353 108 369 142
rect -561 101 369 108
rect 595 142 653 148
rect 595 108 607 142
rect 641 108 653 142
rect 595 102 653 108
rect -695 58 -649 70
rect -695 0 -689 58
rect -701 -7 -689 0
rect -655 0 -649 58
rect -599 58 -553 70
rect -599 0 -593 58
rect -655 -7 -593 0
rect -559 0 -553 58
rect -503 58 -457 70
rect -559 -7 -547 0
rect -701 -63 -699 -7
rect -645 -63 -603 -7
rect -549 -63 -547 -7
rect -701 -70 -547 -63
rect -503 -58 -497 58
rect -463 -58 -457 58
rect -407 58 -361 70
rect -407 0 -401 58
rect -503 -70 -457 -58
rect -413 -7 -401 0
rect -367 0 -361 58
rect -311 58 -265 70
rect -367 -7 -355 0
rect -413 -63 -411 -7
rect -357 -63 -355 -7
rect -413 -70 -355 -63
rect -311 -58 -305 58
rect -271 -58 -265 58
rect -215 58 -169 70
rect -215 0 -209 58
rect -311 -70 -265 -58
rect -221 -7 -209 0
rect -175 0 -169 58
rect -119 58 -73 70
rect -175 -7 -163 0
rect -221 -63 -219 -7
rect -165 -63 -163 -7
rect -221 -70 -163 -63
rect -119 -58 -113 58
rect -79 -58 -73 58
rect -23 58 23 70
rect -23 0 -17 58
rect -119 -70 -73 -58
rect -29 -7 -17 0
rect 17 0 23 58
rect 73 58 119 70
rect 17 -7 29 0
rect -29 -63 -27 -7
rect 27 -63 29 -7
rect -29 -70 29 -63
rect 73 -58 79 58
rect 113 -58 119 58
rect 169 58 215 70
rect 169 0 175 58
rect 73 -70 119 -58
rect 163 -7 175 0
rect 209 0 215 58
rect 265 58 311 70
rect 209 -7 221 0
rect 163 -63 165 -7
rect 219 -63 221 -7
rect 163 -70 221 -63
rect 265 -58 271 58
rect 305 -58 311 58
rect 361 58 407 70
rect 361 0 367 58
rect 265 -70 311 -58
rect 355 -7 367 0
rect 401 0 407 58
rect 457 58 503 70
rect 401 -7 413 0
rect 355 -63 357 -7
rect 411 -63 413 -7
rect 355 -70 413 -63
rect 457 -58 463 58
rect 497 -58 503 58
rect 553 58 599 70
rect 553 0 559 58
rect 457 -70 503 -58
rect 547 -7 559 0
rect 593 0 599 58
rect 649 58 695 70
rect 649 0 655 58
rect 593 -7 655 0
rect 689 0 695 58
rect 689 -7 701 0
rect 547 -63 549 -7
rect 603 -63 645 -7
rect 699 -63 701 -7
rect 547 -70 701 -63
rect -653 -108 -595 -102
rect -653 -142 -641 -108
rect -607 -142 -595 -108
rect -653 -148 -595 -142
rect 403 -108 461 -102
rect 499 -108 557 -102
rect 403 -142 415 -108
rect 449 -142 511 -108
rect 545 -142 557 -108
rect 403 -148 461 -142
rect 499 -148 557 -142
<< via1 >>
rect -699 -58 -689 -7
rect -689 -58 -655 -7
rect -655 -58 -645 -7
rect -699 -63 -645 -58
rect -603 -58 -593 -7
rect -593 -58 -559 -7
rect -559 -58 -549 -7
rect -603 -63 -549 -58
rect -411 -58 -401 -7
rect -401 -58 -367 -7
rect -367 -58 -357 -7
rect -411 -63 -357 -58
rect -219 -58 -209 -7
rect -209 -58 -175 -7
rect -175 -58 -165 -7
rect -219 -63 -165 -58
rect -27 -58 -17 -7
rect -17 -58 17 -7
rect 17 -58 27 -7
rect -27 -63 27 -58
rect 165 -58 175 -7
rect 175 -58 209 -7
rect 209 -58 219 -7
rect 165 -63 219 -58
rect 357 -58 367 -7
rect 367 -58 401 -7
rect 401 -58 411 -7
rect 357 -63 411 -58
rect 549 -58 559 -7
rect 559 -58 593 -7
rect 593 -58 603 -7
rect 549 -63 603 -58
rect 645 -58 655 -7
rect 655 -58 689 -7
rect 689 -58 699 -7
rect 645 -63 699 -58
<< metal2 >>
rect -701 -7 -547 0
rect -701 -63 -699 -7
rect -645 -63 -603 -7
rect -549 -28 -547 -7
rect -413 -7 -355 0
rect -413 -28 -411 -7
rect -549 -63 -411 -28
rect -357 -28 -355 -7
rect -221 -7 -163 0
rect -221 -28 -219 -7
rect -357 -63 -219 -28
rect -165 -28 -163 -7
rect -29 -7 29 0
rect -29 -28 -27 -7
rect -165 -63 -27 -28
rect 27 -28 29 -7
rect 163 -7 221 0
rect 163 -28 165 -7
rect 27 -63 165 -28
rect 219 -63 221 -7
rect -701 -70 221 -63
rect 355 -7 413 0
rect 355 -63 357 -7
rect 411 -28 413 -7
rect 547 -7 701 0
rect 547 -28 549 -7
rect 411 -63 549 -28
rect 603 -63 645 -7
rect 699 -63 701 -7
rect 355 -70 701 -63
<< properties >>
string FIXED_BBOX -786 -227 786 227
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.7 l 0.150 m 1 nf 14 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
