magic
tech sky130A
magscale 1 2
timestamp 1652032815
<< error_p >>
rect -365 151 -307 157
rect -365 117 -353 151
rect -365 111 -307 117
rect 307 -117 365 -111
rect 307 -151 319 -117
rect 307 -157 365 -151
<< nwell >>
rect -743 -289 743 289
<< pmos >>
rect -543 -70 -513 70
rect -447 -70 -417 70
rect -351 -70 -321 70
rect -255 -70 -225 70
rect -159 -70 -129 70
rect -63 -70 -33 70
rect 33 -70 63 70
rect 129 -70 159 70
rect 225 -70 255 70
rect 321 -70 351 70
rect 417 -70 447 70
rect 513 -70 543 70
<< pdiff >>
rect -605 58 -543 70
rect -605 -58 -593 58
rect -559 -58 -543 58
rect -605 -70 -543 -58
rect -513 58 -447 70
rect -513 -58 -497 58
rect -463 -58 -447 58
rect -513 -70 -447 -58
rect -417 58 -351 70
rect -417 -58 -401 58
rect -367 -58 -351 58
rect -417 -70 -351 -58
rect -321 58 -255 70
rect -321 -58 -305 58
rect -271 -58 -255 58
rect -321 -70 -255 -58
rect -225 58 -159 70
rect -225 -58 -209 58
rect -175 -58 -159 58
rect -225 -70 -159 -58
rect -129 58 -63 70
rect -129 -58 -113 58
rect -79 -58 -63 58
rect -129 -70 -63 -58
rect -33 58 33 70
rect -33 -58 -17 58
rect 17 -58 33 58
rect -33 -70 33 -58
rect 63 58 129 70
rect 63 -58 79 58
rect 113 -58 129 58
rect 63 -70 129 -58
rect 159 58 225 70
rect 159 -58 175 58
rect 209 -58 225 58
rect 159 -70 225 -58
rect 255 58 321 70
rect 255 -58 271 58
rect 305 -58 321 58
rect 255 -70 321 -58
rect 351 58 417 70
rect 351 -58 367 58
rect 401 -58 417 58
rect 351 -70 417 -58
rect 447 58 513 70
rect 447 -58 463 58
rect 497 -58 513 58
rect 447 -70 513 -58
rect 543 58 605 70
rect 543 -58 559 58
rect 593 -58 605 58
rect 543 -70 605 -58
<< pdiffc >>
rect -593 -58 -559 58
rect -497 -58 -463 58
rect -401 -58 -367 58
rect -305 -58 -271 58
rect -209 -58 -175 58
rect -113 -58 -79 58
rect -17 -58 17 58
rect 79 -58 113 58
rect 175 -58 209 58
rect 271 -58 305 58
rect 367 -58 401 58
rect 463 -58 497 58
rect 559 -58 593 58
<< nsubdiff >>
rect -707 219 -611 253
rect 611 219 707 253
rect -707 157 -673 219
rect 673 157 707 219
rect -707 -219 -673 -157
rect 673 -219 707 -157
rect -707 -253 -611 -219
rect 611 -253 707 -219
<< nsubdiffcont >>
rect -611 219 611 253
rect -707 -157 -673 157
rect 673 -157 707 157
rect -611 -253 611 -219
<< poly >>
rect -369 151 -303 167
rect -177 151 -111 167
rect 399 151 465 167
rect -369 117 -353 151
rect -319 117 -303 151
rect -369 101 -303 117
rect -255 117 -161 151
rect -127 117 -33 151
rect -543 70 -513 96
rect -447 70 -417 96
rect -351 70 -321 101
rect -255 70 -225 117
rect -177 101 -111 117
rect -159 70 -129 101
rect -63 70 -33 117
rect 399 117 415 151
rect 449 117 465 151
rect 399 101 465 117
rect 33 70 63 96
rect 129 70 159 96
rect 225 70 255 96
rect 321 70 351 96
rect 417 70 447 101
rect 513 70 543 96
rect -543 -96 -513 -70
rect -447 -101 -417 -70
rect -351 -96 -321 -70
rect -255 -96 -225 -70
rect -159 -96 -129 -70
rect -63 -96 -33 -70
rect -465 -117 -399 -101
rect -465 -151 -449 -117
rect -415 -151 -399 -117
rect 33 -117 63 -70
rect 129 -101 159 -70
rect 111 -117 177 -101
rect 225 -117 255 -70
rect 321 -101 351 -70
rect 417 -96 447 -70
rect 513 -96 543 -70
rect 33 -151 127 -117
rect 161 -151 255 -117
rect 303 -117 369 -101
rect 303 -151 319 -117
rect 353 -151 369 -117
rect -465 -167 -399 -151
rect 111 -167 177 -151
rect 303 -167 369 -151
<< polycont >>
rect -353 117 -319 151
rect -161 117 -127 151
rect 415 117 449 151
rect -449 -151 -415 -117
rect 127 -151 161 -117
rect 319 -151 353 -117
<< locali >>
rect -707 219 -611 253
rect 611 219 707 253
rect -707 157 -673 219
rect 673 157 707 219
rect -369 117 -353 151
rect -319 117 -303 151
rect -177 117 -161 151
rect -127 117 -111 151
rect 399 117 415 151
rect 449 117 465 151
rect -593 58 -559 74
rect -593 -74 -559 -58
rect -497 58 -463 74
rect -497 -74 -463 -58
rect -401 58 -367 74
rect -401 -74 -367 -58
rect -305 58 -271 74
rect -305 -74 -271 -58
rect -209 58 -175 74
rect -209 -74 -175 -58
rect -113 58 -79 74
rect -113 -74 -79 -58
rect -17 58 17 74
rect -17 -74 17 -58
rect 79 58 113 74
rect 79 -74 113 -58
rect 175 58 209 74
rect 175 -74 209 -58
rect 271 58 305 74
rect 271 -74 305 -58
rect 367 58 401 74
rect 367 -74 401 -58
rect 463 58 497 74
rect 463 -74 497 -58
rect 559 58 593 74
rect 559 -74 593 -58
rect -465 -151 -449 -117
rect -415 -151 -399 -117
rect 111 -151 127 -117
rect 161 -151 177 -117
rect 303 -151 319 -117
rect 353 -151 369 -117
rect -707 -219 -673 -157
rect 673 -219 707 -157
rect -707 -253 -611 -219
rect 611 -253 707 -219
<< viali >>
rect -353 117 -319 151
rect -161 117 -127 151
rect 415 117 449 151
rect -593 -58 -559 58
rect -497 -58 -463 58
rect -401 -58 -367 58
rect -305 -58 -271 58
rect -209 -58 -175 58
rect -113 -58 -79 58
rect -17 -58 17 58
rect 79 -58 113 58
rect 175 -58 209 58
rect 271 -58 305 58
rect 367 -58 401 58
rect 463 -58 497 58
rect 559 -58 593 58
rect -449 -151 -415 -117
rect 127 -151 161 -117
rect 319 -151 353 -117
<< metal1 >>
rect -365 151 -307 157
rect -365 117 -353 151
rect -319 117 -307 151
rect -365 111 -307 117
rect -173 151 -115 157
rect 403 151 461 157
rect -173 117 -161 151
rect -127 117 415 151
rect 449 117 497 151
rect -173 111 -115 117
rect 79 70 113 117
rect 271 70 305 117
rect 403 111 497 117
rect 463 70 497 111
rect -599 58 -553 70
rect -599 -58 -593 58
rect -559 -58 -553 58
rect -599 -70 -553 -58
rect -503 58 -457 70
rect -503 -58 -497 58
rect -463 -58 -457 58
rect -503 -70 -457 -58
rect -417 63 -351 70
rect -417 -63 -407 63
rect -355 -63 -351 63
rect -417 -70 -351 -63
rect -311 58 -265 70
rect -311 -58 -305 58
rect -271 -58 -265 58
rect -311 -70 -265 -58
rect -225 63 -159 70
rect -225 -63 -215 63
rect -163 -63 -159 63
rect -225 -70 -159 -63
rect -119 58 -73 70
rect -119 -58 -113 58
rect -79 -58 -73 58
rect -119 -70 -73 -58
rect -33 63 33 70
rect -33 -63 -23 63
rect 29 -63 33 63
rect -33 -70 33 -63
rect 73 58 119 70
rect 73 -58 79 58
rect 113 -58 119 58
rect 73 -70 119 -58
rect 159 63 225 70
rect 159 -63 169 63
rect 221 -63 225 63
rect 159 -70 225 -63
rect 265 58 311 70
rect 265 -58 271 58
rect 305 -58 311 58
rect 265 -70 311 -58
rect 351 63 417 70
rect 351 -63 361 63
rect 413 -63 417 63
rect 351 -70 417 -63
rect 457 58 503 70
rect 457 -58 463 58
rect 497 -58 503 58
rect 457 -70 503 -58
rect 553 58 599 70
rect 553 -58 559 58
rect 593 -58 599 58
rect 553 -70 599 -58
rect -497 -111 -463 -70
rect -497 -117 -403 -111
rect -305 -117 -271 -70
rect -113 -117 -79 -70
rect 115 -117 173 -111
rect -497 -151 -449 -117
rect -415 -151 127 -117
rect 161 -151 173 -117
rect -461 -157 -403 -151
rect -113 -289 -79 -151
rect 115 -157 173 -151
rect 307 -117 365 -111
rect 307 -151 319 -117
rect 353 -151 365 -117
rect 307 -157 365 -151
rect 463 -185 497 -70
rect 79 -219 497 -185
rect 79 -289 113 -219
<< via1 >>
rect -407 58 -355 63
rect -407 -58 -401 58
rect -401 -58 -367 58
rect -367 -58 -355 58
rect -407 -63 -355 -58
rect -215 58 -163 63
rect -215 -58 -209 58
rect -209 -58 -175 58
rect -175 -58 -163 58
rect -215 -63 -163 -58
rect -23 58 29 63
rect -23 -58 -17 58
rect -17 -58 17 58
rect 17 -58 29 58
rect -23 -63 29 -58
rect 169 58 221 63
rect 169 -58 175 58
rect 175 -58 209 58
rect 209 -58 221 58
rect 169 -63 221 -58
rect 361 58 413 63
rect 361 -58 367 58
rect 367 -58 401 58
rect 401 -58 413 58
rect 361 -63 413 -58
<< metal2 >>
rect -417 63 -351 70
rect -417 17 -407 63
rect -661 -17 -407 17
rect -417 -63 -407 -17
rect -355 17 -351 63
rect -225 63 -159 70
rect -225 17 -215 63
rect -355 -17 -215 17
rect -355 -63 -351 -17
rect -417 -70 -351 -63
rect -225 -63 -215 -17
rect -163 17 -159 63
rect -33 63 33 70
rect -33 17 -23 63
rect -163 -17 -23 17
rect -163 -63 -159 -17
rect -225 -70 -159 -63
rect -33 -63 -23 -17
rect 29 17 33 63
rect 159 63 225 70
rect 159 17 169 63
rect 29 -17 169 17
rect 29 -63 33 -17
rect -33 -70 33 -63
rect 159 -63 169 -17
rect 221 17 225 63
rect 351 63 417 70
rect 351 17 361 63
rect 221 -17 361 17
rect 221 -63 225 -17
rect 159 -70 225 -63
rect 351 -63 361 -17
rect 413 -63 417 63
rect 351 -70 417 -63
<< properties >>
string FIXED_BBOX -690 -236 690 236
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.7 l 0.15 m 1 nf 12 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
