magic
tech sky130A
magscale 1 2
timestamp 1660307144
<< nwell >>
rect 1786 261 1862 582
<< locali >>
rect 18 -1755 84 -1735
rect 18 -1789 32 -1755
rect 66 -1789 84 -1755
rect 18 -1803 84 -1789
<< viali >>
rect 32 215 66 249
rect 289 221 323 255
rect 1928 220 1962 254
rect 1396 130 1430 164
rect 2020 85 2054 255
rect 2112 221 2146 255
rect 32 -453 66 -419
rect 289 -447 323 -413
rect 1396 -538 1430 -504
rect 32 -1121 66 -1087
rect 289 -1115 323 -1081
rect 1396 -1206 1430 -1172
rect 1679 -1695 1713 -1661
rect 32 -1789 66 -1755
rect 289 -1789 323 -1755
rect 1396 -1874 1430 -1840
<< metal1 >>
rect 14 570 78 576
rect 14 518 20 570
rect 72 518 78 570
rect 1748 520 1900 568
rect 14 512 78 518
rect 1025 289 2058 331
rect -114 255 -108 258
rect -127 209 -108 255
rect -114 206 -108 209
rect -56 255 -50 258
rect 22 255 76 261
rect -56 249 76 255
rect -56 215 32 249
rect 66 215 76 249
rect -56 209 76 215
rect 274 255 335 264
rect 274 221 289 255
rect 323 253 335 255
rect 1025 253 1067 289
rect 2008 267 2058 289
rect 323 221 1067 253
rect 274 211 1067 221
rect 1804 254 1979 260
rect 1804 220 1928 254
rect 1962 220 1979 254
rect 1804 216 1979 220
rect -56 206 -50 209
rect -105 198 -59 206
rect 22 203 76 209
rect 1381 173 1445 179
rect 1381 121 1387 173
rect 1439 121 1445 173
rect 1381 115 1445 121
rect 14 -98 78 -92
rect 14 -150 20 -98
rect 72 -150 78 -98
rect 14 -156 78 -150
rect -105 -410 -59 -408
rect -114 -462 -108 -410
rect -56 -413 -50 -410
rect 22 -413 76 -407
rect -56 -419 76 -413
rect -56 -453 32 -419
rect 66 -453 76 -419
rect -56 -459 76 -453
rect -56 -462 -50 -459
rect -105 -474 -59 -462
rect 22 -465 76 -459
rect 274 -410 338 -404
rect 274 -462 280 -410
rect 332 -462 338 -410
rect 274 -468 338 -462
rect 274 -513 320 -468
rect 1804 -489 1848 216
rect 1919 211 1979 216
rect 2008 255 2066 267
rect 2008 85 2020 255
rect 2054 85 2066 255
rect 2095 260 2155 264
rect 2095 255 2279 260
rect 2095 221 2112 255
rect 2146 221 2279 255
rect 2095 216 2279 221
rect 2095 211 2155 216
rect 2008 76 2066 85
rect 1913 26 1977 32
rect 1913 -26 1919 26
rect 1971 -26 1977 26
rect 1913 -32 1977 -26
rect 1387 -495 1848 -489
rect -200 -559 320 -513
rect 1381 -547 1387 -496
rect 1439 -533 1848 -495
rect 1439 -547 1445 -533
rect 1381 -553 1445 -547
rect -200 -1749 -154 -559
rect 14 -766 78 -760
rect 14 -818 20 -766
rect 72 -818 78 -766
rect 14 -824 78 -818
rect -114 -1130 -108 -1078
rect -56 -1081 -50 -1078
rect 22 -1081 76 -1075
rect -56 -1087 76 -1081
rect -56 -1121 32 -1087
rect 66 -1121 76 -1087
rect -56 -1127 76 -1121
rect -56 -1130 -50 -1127
rect 22 -1133 76 -1127
rect 274 -1078 338 -1072
rect 274 -1130 280 -1078
rect 332 -1130 338 -1078
rect 274 -1136 338 -1130
rect 2235 -1157 2279 216
rect 1381 -1172 2279 -1157
rect 1381 -1206 1396 -1172
rect 1430 -1201 2279 -1172
rect 1430 -1206 1445 -1201
rect 1381 -1221 1445 -1206
rect 1670 -1310 1734 -1304
rect 1670 -1362 1676 -1310
rect 1728 -1362 1734 -1310
rect 1670 -1368 1734 -1362
rect 14 -1434 78 -1428
rect 14 -1486 20 -1434
rect 72 -1486 78 -1434
rect 14 -1492 78 -1486
rect 1669 -1661 1723 -1649
rect 1669 -1695 1679 -1661
rect 1713 -1695 1723 -1661
rect 1669 -1707 1723 -1695
rect 22 -1749 76 -1743
rect -200 -1755 76 -1749
rect -200 -1789 32 -1755
rect 66 -1789 76 -1755
rect -200 -1795 76 -1789
rect 22 -1801 76 -1795
rect 279 -1749 333 -1743
rect 1673 -1749 1719 -1707
rect 279 -1755 1719 -1749
rect 279 -1789 289 -1755
rect 323 -1789 1719 -1755
rect 279 -1794 1719 -1789
rect 279 -1795 1718 -1794
rect 279 -1801 333 -1795
rect 1386 -1834 1440 -1828
rect 1386 -1840 1925 -1834
rect 1386 -1874 1396 -1840
rect 1430 -1874 1925 -1840
rect 1386 -1880 1925 -1874
rect 1386 -1886 1440 -1880
<< via1 >>
rect 20 518 72 570
rect -108 206 -56 258
rect 1387 164 1439 173
rect 1387 130 1396 164
rect 1396 130 1430 164
rect 1430 130 1439 164
rect 1387 121 1439 130
rect 1676 -26 1728 26
rect 20 -150 72 -98
rect -108 -462 -56 -410
rect 280 -413 332 -410
rect 280 -447 289 -413
rect 289 -447 323 -413
rect 323 -447 332 -413
rect 280 -462 332 -447
rect 1919 -26 1971 26
rect 1387 -504 1439 -495
rect 1387 -538 1396 -504
rect 1396 -538 1430 -504
rect 1430 -538 1439 -504
rect 1387 -547 1439 -538
rect 1676 -694 1728 -642
rect 20 -818 72 -766
rect -108 -1130 -56 -1078
rect 280 -1081 332 -1078
rect 280 -1115 289 -1081
rect 289 -1115 323 -1081
rect 323 -1115 332 -1081
rect 280 -1130 332 -1115
rect 1676 -1362 1728 -1310
rect 20 -1486 72 -1434
rect 1676 -2030 1728 -1978
<< metal2 >>
rect 22 576 70 694
rect 14 570 78 576
rect 14 518 20 570
rect 72 518 78 570
rect 14 512 78 518
rect -108 258 -56 264
rect -108 200 -56 206
rect -105 -404 -59 200
rect 22 -92 70 512
rect 1381 173 1445 179
rect 1381 121 1387 173
rect 1439 121 1445 173
rect 1381 115 1445 121
rect 1381 88 1437 115
rect 282 40 1437 88
rect 14 -98 78 -92
rect 14 -150 20 -98
rect 72 -150 78 -98
rect 14 -156 78 -150
rect -108 -410 -56 -404
rect -108 -468 -56 -462
rect -105 -1072 -59 -468
rect 22 -760 70 -156
rect 282 -404 330 40
rect 1678 32 1726 694
rect 1670 26 1734 32
rect 1670 -26 1676 26
rect 1728 25 1734 26
rect 1913 26 1977 32
rect 1728 24 1781 25
rect 1913 24 1919 26
rect 1728 -23 1919 24
rect 1728 -26 1734 -23
rect 1781 -24 1919 -23
rect 1670 -32 1734 -26
rect 1913 -26 1919 -24
rect 1971 -26 1977 26
rect 1913 -32 1977 -26
rect 274 -410 338 -404
rect 274 -462 280 -410
rect 332 -462 338 -410
rect 274 -468 338 -462
rect 1381 -495 1445 -489
rect 1381 -547 1387 -495
rect 1439 -547 1445 -495
rect 1381 -553 1445 -547
rect 1381 -580 1437 -553
rect 282 -628 1437 -580
rect 14 -766 78 -760
rect 14 -818 20 -766
rect 72 -818 78 -766
rect 14 -824 78 -818
rect -108 -1078 -56 -1072
rect -108 -1136 -56 -1130
rect 22 -1428 70 -824
rect 282 -1072 330 -628
rect 1678 -636 1726 -32
rect 1670 -642 1734 -636
rect 1670 -694 1676 -642
rect 1728 -694 1734 -642
rect 1670 -700 1734 -694
rect 274 -1078 338 -1072
rect 274 -1130 280 -1078
rect 332 -1130 338 -1078
rect 274 -1136 338 -1130
rect 1678 -1304 1726 -700
rect 1670 -1310 1734 -1304
rect 1670 -1362 1676 -1310
rect 1728 -1362 1734 -1310
rect 1670 -1368 1734 -1362
rect 14 -1434 78 -1428
rect 14 -1486 20 -1434
rect 72 -1486 78 -1434
rect 14 -1492 78 -1486
rect 1678 -1972 1726 -1368
rect 1670 -1978 1734 -1972
rect 1670 -2030 1676 -1978
rect 1728 -2030 1734 -1978
rect 1670 -2036 1734 -2030
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_0 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 0 0 1 0
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_1
timestamp 1644511149
transform 1 0 0 0 1 -668
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_2
timestamp 1644511149
transform 1 0 0 0 1 -1336
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_3
timestamp 1644511149
transform 1 0 0 0 1 -2004
box -38 -48 1786 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_0 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1900 0 1 0
box -38 -48 314 592
<< labels >>
rlabel metal1 -127 209 -51 255 0 clkin
rlabel metal2 22 650 70 694 0 VPWR
rlabel metal2 1678 650 1726 694 6 VGND
rlabel metal1 -105 -1795 -61 -1749 5 s1
rlabel metal1 1881 -1880 1925 -1834 5 s2
<< end >>
