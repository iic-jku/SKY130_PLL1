magic
tech sky130A
magscale 1 2
timestamp 1668357910
<< pwell >>
rect -743 -280 743 280
<< nmos >>
rect -543 -70 -513 70
rect -447 -70 -417 70
rect -351 -70 -321 70
rect -255 -70 -225 70
rect -159 -70 -129 70
rect -63 -70 -33 70
rect 33 -70 63 70
rect 129 -70 159 70
rect 225 -70 255 70
rect 321 -70 351 70
rect 417 -70 447 70
rect 513 -70 543 70
<< ndiff >>
rect -605 58 -543 70
rect -605 -58 -593 58
rect -559 -58 -543 58
rect -605 -70 -543 -58
rect -513 58 -447 70
rect -513 -58 -497 58
rect -463 -58 -447 58
rect -513 -70 -447 -58
rect -417 58 -351 70
rect -417 -58 -401 58
rect -367 -58 -351 58
rect -417 -70 -351 -58
rect -321 58 -255 70
rect -321 -58 -305 58
rect -271 -58 -255 58
rect -321 -70 -255 -58
rect -225 58 -159 70
rect -225 -58 -209 58
rect -175 -58 -159 58
rect -225 -70 -159 -58
rect -129 58 -63 70
rect -129 -58 -113 58
rect -79 -58 -63 58
rect -129 -70 -63 -58
rect -33 58 33 70
rect -33 -58 -17 58
rect 17 -58 33 58
rect -33 -70 33 -58
rect 63 58 129 70
rect 63 -58 79 58
rect 113 -58 129 58
rect 63 -70 129 -58
rect 159 58 225 70
rect 159 -58 175 58
rect 209 -58 225 58
rect 159 -70 225 -58
rect 255 58 321 70
rect 255 -58 271 58
rect 305 -58 321 58
rect 255 -70 321 -58
rect 351 58 417 70
rect 351 -58 367 58
rect 401 -58 417 58
rect 351 -70 417 -58
rect 447 58 513 70
rect 447 -58 463 58
rect 497 -58 513 58
rect 447 -70 513 -58
rect 543 58 605 70
rect 543 -58 559 58
rect 593 -58 605 58
rect 543 -70 605 -58
<< ndiffc >>
rect -593 -58 -559 58
rect -497 -58 -463 58
rect -401 -58 -367 58
rect -305 -58 -271 58
rect -209 -58 -175 58
rect -113 -58 -79 58
rect -17 -58 17 58
rect 79 -58 113 58
rect 175 -58 209 58
rect 271 -58 305 58
rect 367 -58 401 58
rect 463 -58 497 58
rect 559 -58 593 58
<< psubdiff >>
rect -707 210 -611 244
rect 611 210 707 244
rect -707 148 -673 210
rect 673 148 707 210
rect -707 -210 -673 -148
rect 673 -210 707 -148
rect -707 -244 -611 -210
rect 611 -244 707 -210
<< psubdiffcont >>
rect -611 210 611 244
rect -707 -148 -673 148
rect 673 -148 707 148
rect -611 -244 611 -210
<< poly >>
rect -465 142 465 158
rect -465 108 -449 142
rect -415 108 -353 142
rect -319 108 -257 142
rect -223 108 -161 142
rect -127 108 -65 142
rect -31 108 31 142
rect 65 108 127 142
rect 161 108 223 142
rect 257 108 319 142
rect 353 108 415 142
rect 449 108 465 142
rect -543 70 -513 96
rect -465 92 465 108
rect -447 70 -417 92
rect -351 70 -321 92
rect -255 70 -225 92
rect -159 70 -129 92
rect -63 70 -33 92
rect 33 70 63 92
rect 129 70 159 92
rect 225 70 255 92
rect 321 70 351 92
rect 417 70 447 92
rect 513 70 543 96
rect -543 -92 -513 -70
rect -561 -108 -495 -92
rect -447 -96 -417 -70
rect -351 -96 -321 -70
rect -255 -96 -225 -70
rect -159 -97 -129 -70
rect -63 -96 -33 -70
rect 33 -96 63 -70
rect 129 -96 159 -70
rect 225 -96 255 -70
rect 321 -96 351 -70
rect 417 -96 447 -70
rect 513 -92 543 -70
rect -561 -142 -545 -108
rect -511 -142 -495 -108
rect -561 -158 -495 -142
rect 495 -108 561 -92
rect 495 -142 511 -108
rect 545 -142 561 -108
rect 495 -158 561 -142
<< polycont >>
rect -449 108 -415 142
rect -353 108 -319 142
rect -257 108 -223 142
rect -161 108 -127 142
rect -65 108 -31 142
rect 31 108 65 142
rect 127 108 161 142
rect 223 108 257 142
rect 319 108 353 142
rect 415 108 449 142
rect -545 -142 -511 -108
rect 511 -142 545 -108
<< locali >>
rect -707 210 -611 244
rect 611 210 707 244
rect -707 148 -673 210
rect 673 148 707 210
rect -465 108 -449 142
rect -415 108 -353 142
rect -319 108 -257 142
rect -223 108 -161 142
rect -127 108 -65 142
rect -31 108 31 142
rect 65 108 127 142
rect 161 108 223 142
rect 257 108 319 142
rect 353 108 415 142
rect 449 108 465 142
rect -707 -210 -673 -148
rect -593 58 -559 74
rect -593 -108 -559 -58
rect -497 58 -463 74
rect -497 -74 -463 -58
rect -401 58 -367 74
rect -401 -74 -367 -58
rect -305 58 -271 74
rect -305 -74 -271 -58
rect -209 58 -175 74
rect -209 -74 -175 -58
rect -113 58 -79 74
rect -113 -74 -79 -58
rect -17 58 17 74
rect -17 -74 17 -58
rect 79 58 113 74
rect 79 -74 113 -58
rect 175 58 209 74
rect 175 -74 209 -58
rect 271 58 305 74
rect 271 -74 305 -58
rect 367 58 401 74
rect 367 -74 401 -58
rect 463 58 497 74
rect 463 -74 497 -58
rect 559 58 593 74
rect 559 -108 593 -58
rect -593 -142 -545 -108
rect -511 -142 -495 -108
rect 495 -142 511 -108
rect 545 -142 593 -108
rect -593 -210 -559 -142
rect 559 -210 593 -142
rect 673 -210 707 -148
rect -707 -244 -611 -210
rect 611 -244 707 -210
<< viali >>
rect -449 108 -415 142
rect -353 108 -319 142
rect -257 108 -223 142
rect -161 108 -127 142
rect -65 108 -31 142
rect 31 108 65 142
rect 127 108 161 142
rect 223 108 257 142
rect 319 108 353 142
rect 415 108 449 142
rect -593 -58 -559 58
rect -497 -58 -463 58
rect -401 -58 -367 58
rect -305 -58 -271 58
rect -209 -58 -175 58
rect -113 -58 -79 58
rect -17 -58 17 58
rect 79 -58 113 58
rect 175 -58 209 58
rect 271 -58 305 58
rect 367 -58 401 58
rect 463 -58 497 58
rect 559 -58 593 58
rect -545 -142 -511 -108
rect 511 -142 545 -108
<< metal1 >>
rect -461 142 -403 148
rect -365 142 -307 148
rect -269 142 -211 148
rect -173 142 -115 148
rect -77 142 -19 148
rect 19 142 77 148
rect 115 142 173 148
rect 211 142 269 148
rect 307 142 365 148
rect 403 142 461 148
rect -465 108 -449 142
rect -415 108 -353 142
rect -319 108 -257 142
rect -223 108 -161 142
rect -127 108 -65 142
rect -31 108 31 142
rect 65 108 127 142
rect 161 108 223 142
rect 257 108 319 142
rect 353 108 415 142
rect 449 108 465 142
rect -461 102 -403 108
rect -365 102 -307 108
rect -269 102 -211 108
rect -173 102 -115 108
rect -77 102 -19 108
rect 19 102 77 108
rect 115 102 173 108
rect 211 102 269 108
rect 307 102 365 108
rect 403 102 461 108
rect -599 58 -553 70
rect -599 0 -593 58
rect -604 -7 -593 0
rect -559 0 -553 58
rect -503 58 -457 70
rect -503 0 -497 58
rect -559 -7 -497 0
rect -463 0 -457 58
rect -407 58 -361 70
rect -463 -7 -452 0
rect -604 -63 -603 -7
rect -550 -63 -507 -7
rect -454 -63 -452 -7
rect -604 -70 -452 -63
rect -407 -58 -401 58
rect -367 -58 -361 58
rect -311 58 -265 70
rect -311 0 -305 58
rect -407 -70 -361 -58
rect -316 -7 -305 0
rect -271 0 -265 58
rect -215 58 -169 70
rect -271 -7 -260 0
rect -316 -63 -315 -7
rect -262 -63 -260 -7
rect -316 -70 -260 -63
rect -215 -58 -209 58
rect -175 -58 -169 58
rect -119 58 -73 70
rect -119 0 -113 58
rect -215 -70 -169 -58
rect -124 -7 -113 0
rect -79 0 -73 58
rect -23 58 23 70
rect -79 -7 -68 0
rect -124 -63 -123 -7
rect -70 -63 -68 -7
rect -124 -70 -68 -63
rect -23 -58 -17 58
rect 17 -58 23 58
rect 73 58 119 70
rect 73 0 79 58
rect -23 -70 23 -58
rect 68 -7 79 0
rect 113 0 119 58
rect 169 58 215 70
rect 113 -7 124 0
rect 68 -63 69 -7
rect 122 -63 124 -7
rect 68 -70 124 -63
rect 169 -58 175 58
rect 209 -58 215 58
rect 265 58 311 70
rect 265 0 271 58
rect 169 -70 215 -58
rect 260 -7 271 0
rect 305 0 311 58
rect 361 58 407 70
rect 305 -7 316 0
rect 260 -63 261 -7
rect 314 -63 316 -7
rect 260 -70 316 -63
rect 361 -58 367 58
rect 401 -58 407 58
rect 457 58 503 70
rect 457 0 463 58
rect 361 -70 407 -58
rect 452 -7 463 0
rect 497 0 503 58
rect 553 58 599 70
rect 553 0 559 58
rect 497 -7 559 0
rect 593 0 599 58
rect 593 -7 604 0
rect 452 -63 453 -7
rect 506 -63 549 -7
rect 602 -63 604 -7
rect 452 -70 604 -63
rect -593 -102 -557 -70
rect 557 -102 593 -70
rect -593 -108 -499 -102
rect -593 -142 -545 -108
rect -511 -142 -499 -108
rect -593 -148 -499 -142
rect 499 -108 593 -102
rect 499 -142 511 -108
rect 545 -142 593 -108
rect 499 -148 593 -142
<< via1 >>
rect -603 -58 -593 -7
rect -593 -58 -559 -7
rect -559 -58 -550 -7
rect -603 -63 -550 -58
rect -507 -58 -497 -7
rect -497 -58 -463 -7
rect -463 -58 -454 -7
rect -507 -63 -454 -58
rect -315 -58 -305 -7
rect -305 -58 -271 -7
rect -271 -58 -262 -7
rect -315 -63 -262 -58
rect -123 -58 -113 -7
rect -113 -58 -79 -7
rect -79 -58 -70 -7
rect -123 -63 -70 -58
rect 69 -58 79 -7
rect 79 -58 113 -7
rect 113 -58 122 -7
rect 69 -63 122 -58
rect 261 -58 271 -7
rect 271 -58 305 -7
rect 305 -58 314 -7
rect 261 -63 314 -58
rect 453 -58 463 -7
rect 463 -58 497 -7
rect 497 -58 506 -7
rect 453 -63 506 -58
rect 549 -58 559 -7
rect 559 -58 593 -7
rect 593 -58 602 -7
rect 549 -63 602 -58
<< metal2 >>
rect -604 -7 -452 0
rect -604 -63 -603 -7
rect -550 -63 -507 -7
rect -454 -28 -452 -7
rect -316 -7 -260 0
rect -316 -28 -315 -7
rect -454 -63 -315 -28
rect -262 -28 -260 -7
rect -124 -7 -68 0
rect -124 -28 -123 -7
rect -262 -63 -123 -28
rect -70 -28 -68 -7
rect 68 -7 124 0
rect 68 -28 69 -7
rect -70 -63 69 -28
rect 122 -28 124 -7
rect 260 -7 316 0
rect 260 -28 261 -7
rect 122 -63 261 -28
rect 314 -28 316 -7
rect 452 -7 604 0
rect 452 -28 453 -7
rect 314 -63 453 -28
rect 506 -63 549 -7
rect 602 -63 604 -7
rect -604 -70 604 -63
<< properties >>
string FIXED_BBOX -690 -227 690 227
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.7 l 0.150 m 1 nf 12 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
