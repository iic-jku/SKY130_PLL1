magic
tech sky130A
magscale 1 2
timestamp 1666520455
<< metal1 >>
rect 70 2104 186 2138
rect 724 2104 1096 2138
rect 1634 2104 2006 2138
rect 70 1885 104 2104
rect -139 1879 631 1885
rect -139 1827 573 1879
rect 625 1827 631 1879
rect -139 1821 631 1827
rect -139 1462 -75 1821
rect -139 1392 -75 1398
rect -42 1677 952 1719
rect -42 539 0 1677
rect 1788 1672 1794 1724
rect 1846 1672 1852 1724
rect 423 1517 429 1569
rect 481 1560 487 1569
rect 481 1526 570 1560
rect 481 1517 487 1526
rect 2730 1406 2788 1412
rect 1897 1310 1903 1319
rect 820 1276 1192 1310
rect 1538 1276 1903 1310
rect 1897 1267 1903 1276
rect 1955 1310 1961 1319
rect 1955 1276 2102 1310
rect 1955 1267 1961 1276
rect 2730 1000 2788 1348
rect 724 966 1096 1000
rect 1634 966 2006 1000
rect 2544 966 2788 1000
rect 878 534 884 586
rect 936 534 942 586
rect 1788 534 1794 586
rect 1846 534 1852 586
rect 963 393 1015 399
rect 963 335 1015 341
rect 1873 388 1925 394
rect 972 172 1006 335
rect 1873 330 1925 336
rect 1882 172 1916 330
rect 2730 268 2788 966
rect 2730 204 2788 210
rect 628 138 1192 172
rect 1538 138 2102 172
<< via1 >>
rect 573 1827 625 1879
rect -139 1398 -75 1462
rect 1794 1672 1846 1724
rect 429 1517 481 1569
rect 2730 1348 2788 1406
rect 1903 1267 1955 1319
rect 884 534 936 586
rect 1794 534 1846 586
rect 963 341 1015 393
rect 1873 336 1925 388
rect 2730 210 2788 268
<< metal2 >>
rect 772 1987 1048 2057
rect 426 1571 484 1917
rect 567 1879 676 1882
rect 567 1827 573 1879
rect 625 1827 676 1879
rect 567 1824 676 1827
rect -139 1569 484 1571
rect -139 1517 429 1569
rect 481 1517 484 1569
rect -139 1513 484 1517
rect -145 1398 -139 1462
rect -75 1398 -69 1462
rect -139 268 -75 1398
rect 80 861 138 1513
rect 429 1511 481 1513
rect 618 1488 676 1824
rect 1794 1724 1846 1730
rect 1788 1677 1794 1719
rect 1794 1666 1846 1672
rect 868 1348 1144 1418
rect 1900 1319 1958 2057
rect 2592 1999 2794 2057
rect 2730 1677 2772 1719
rect 2496 1348 2730 1406
rect 2788 1348 2794 1406
rect 1900 1267 1903 1319
rect 1955 1267 1958 1319
rect 1900 919 1958 1267
rect 772 849 1048 919
rect 1682 849 1958 919
rect 884 586 936 592
rect 878 539 884 581
rect 884 528 936 534
rect 972 393 1006 849
rect 1794 586 1846 592
rect 1788 539 1794 581
rect 1794 528 1846 534
rect 957 341 963 393
rect 1015 341 1021 393
rect 1882 388 1916 849
rect 2730 539 2772 581
rect 1867 336 1873 388
rect 1925 336 1931 388
rect -139 210 234 268
rect 676 210 1144 280
rect 1586 210 2054 280
rect 2496 210 2730 268
rect 2788 210 2794 268
use simple_inv  simple_inv_0 /foss/designs/ma2022
timestamp 1660926584
transform 1 0 53 0 1 613
box -53 -613 857 525
use simple_inv  simple_inv_1
timestamp 1660926584
transform 1 0 963 0 1 613
box -53 -613 857 525
use simple_inv  simple_inv_2
timestamp 1660926584
transform 1 0 1873 0 1 613
box -53 -613 857 525
use simple_inv  simple_inv_3
timestamp 1660926584
transform 1 0 1873 0 1 1751
box -53 -613 857 525
use simple_inv  simple_inv_4
timestamp 1660926584
transform 1 0 963 0 1 1751
box -53 -613 857 525
use sinv_n  sinv_n_0 /foss/designs/ma2022
timestamp 1660926584
transform 1 0 647 0 1 1418
box -359 -280 359 280
use sinv_p  sinv_p_0 /foss/designs/ma2022
timestamp 1660926584
transform 1 0 455 0 1 1987
box -455 -289 455 289
<< labels >>
rlabel metal2 2730 539 2772 581 0 nclk
rlabel metal2 2730 1677 2772 1719 0 clk
rlabel metal1 -139 1821 -75 1885 7 vss
rlabel metal2 2736 1999 2794 2057 5 vdd
rlabel metal1 -42 1677 0 1719 6 clk_in
<< end >>
