magic
tech sky130A
magscale 1 2
timestamp 1654967793
<< nwell >>
rect -887 -289 887 289
<< pmos >>
rect -687 -70 -657 70
rect -591 -70 -561 70
rect -495 -70 -465 70
rect -399 -70 -369 70
rect -303 -70 -273 70
rect -207 -70 -177 70
rect -111 -70 -81 70
rect -15 -70 15 70
rect 81 -70 111 70
rect 177 -70 207 70
rect 273 -70 303 70
rect 369 -70 399 70
rect 465 -70 495 70
rect 561 -70 591 70
rect 657 -70 687 70
<< pdiff >>
rect -753 58 -687 70
rect -753 -58 -737 58
rect -703 -58 -687 58
rect -753 -70 -687 -58
rect -657 58 -591 70
rect -657 -58 -641 58
rect -607 -58 -591 58
rect -657 -70 -591 -58
rect -561 58 -495 70
rect -561 -58 -545 58
rect -511 -58 -495 58
rect -561 -70 -495 -58
rect -465 58 -399 70
rect -465 -58 -449 58
rect -415 -58 -399 58
rect -465 -70 -399 -58
rect -369 58 -303 70
rect -369 -58 -353 58
rect -319 -58 -303 58
rect -369 -70 -303 -58
rect -273 58 -207 70
rect -273 -58 -257 58
rect -223 -58 -207 58
rect -273 -70 -207 -58
rect -177 58 -111 70
rect -177 -58 -161 58
rect -127 -58 -111 58
rect -177 -70 -111 -58
rect -81 58 -15 70
rect -81 -58 -65 58
rect -31 -58 -15 58
rect -81 -70 -15 -58
rect 15 58 81 70
rect 15 -58 31 58
rect 65 -58 81 58
rect 15 -70 81 -58
rect 111 58 177 70
rect 111 -58 127 58
rect 161 -58 177 58
rect 111 -70 177 -58
rect 207 58 273 70
rect 207 -58 223 58
rect 257 -58 273 58
rect 207 -70 273 -58
rect 303 58 369 70
rect 303 -58 319 58
rect 353 -58 369 58
rect 303 -70 369 -58
rect 399 58 465 70
rect 399 -58 415 58
rect 449 -58 465 58
rect 399 -70 465 -58
rect 495 58 561 70
rect 495 -58 511 58
rect 545 -58 561 58
rect 495 -70 561 -58
rect 591 58 657 70
rect 591 -58 607 58
rect 641 -58 657 58
rect 591 -70 657 -58
rect 687 58 753 70
rect 687 -58 703 58
rect 737 -58 753 58
rect 687 -70 753 -58
<< pdiffc >>
rect -737 -58 -703 58
rect -641 -58 -607 58
rect -545 -58 -511 58
rect -449 -58 -415 58
rect -353 -58 -319 58
rect -257 -58 -223 58
rect -161 -58 -127 58
rect -65 -58 -31 58
rect 31 -58 65 58
rect 127 -58 161 58
rect 223 -58 257 58
rect 319 -58 353 58
rect 415 -58 449 58
rect 511 -58 545 58
rect 607 -58 641 58
rect 703 -58 737 58
<< nsubdiff >>
rect -851 219 -755 253
rect 755 219 851 253
rect -851 157 -817 219
rect 817 157 851 219
rect -851 -219 -817 -157
rect 817 -219 851 -157
rect -851 -253 -755 -219
rect 755 -253 851 -219
<< nsubdiffcont >>
rect -755 219 755 253
rect -851 -157 -817 157
rect 817 -157 851 157
rect -755 -253 755 -219
<< poly >>
rect -609 151 609 167
rect -609 117 -593 151
rect -559 117 -497 151
rect -463 117 -401 151
rect -367 117 -305 151
rect -271 117 -209 151
rect -175 117 -113 151
rect -79 117 -17 151
rect 17 117 79 151
rect 113 117 175 151
rect 209 117 271 151
rect 305 117 367 151
rect 401 117 463 151
rect 497 117 559 151
rect 593 117 609 151
rect -609 101 609 117
rect -687 70 -657 96
rect -591 70 -561 101
rect -495 70 -465 101
rect -399 70 -369 101
rect -303 70 -273 101
rect -207 70 -177 101
rect -111 70 -81 101
rect -15 70 15 101
rect 81 70 111 101
rect 177 70 207 101
rect 273 70 303 101
rect 369 70 399 101
rect 465 70 495 101
rect 561 70 591 101
rect 657 70 687 96
rect -687 -101 -657 -70
rect -591 -96 -561 -70
rect -495 -96 -465 -70
rect -399 -96 -369 -70
rect -303 -96 -273 -70
rect -207 -96 -177 -70
rect -111 -96 -81 -70
rect -15 -96 15 -70
rect 81 -96 111 -70
rect 177 -96 207 -70
rect 273 -96 303 -70
rect 369 -96 399 -70
rect 465 -96 495 -70
rect 561 -96 591 -70
rect 657 -101 687 -70
rect -705 -117 -639 -101
rect -705 -151 -689 -117
rect -655 -151 -639 -117
rect -705 -167 -639 -151
rect 639 -117 705 -101
rect 639 -151 655 -117
rect 689 -151 705 -117
rect 639 -167 705 -151
<< polycont >>
rect -593 117 -559 151
rect -497 117 -463 151
rect -401 117 -367 151
rect -305 117 -271 151
rect -209 117 -175 151
rect -113 117 -79 151
rect -17 117 17 151
rect 79 117 113 151
rect 175 117 209 151
rect 271 117 305 151
rect 367 117 401 151
rect 463 117 497 151
rect 559 117 593 151
rect -689 -151 -655 -117
rect 655 -151 689 -117
<< locali >>
rect -851 219 -755 253
rect 755 219 851 253
rect -851 157 -817 219
rect 817 157 851 219
rect -609 117 -593 151
rect -559 117 -497 151
rect -463 117 -401 151
rect -367 117 -305 151
rect -271 117 -209 151
rect -175 117 -113 151
rect -79 117 -17 151
rect 17 117 79 151
rect 113 117 175 151
rect 209 117 271 151
rect 305 117 367 151
rect 401 117 463 151
rect 497 117 559 151
rect 593 117 609 151
rect -737 58 -703 74
rect -737 -74 -703 -58
rect -641 58 -607 74
rect -641 -74 -607 -58
rect -545 58 -511 74
rect -545 -74 -511 -58
rect -449 58 -415 74
rect -449 -74 -415 -58
rect -353 58 -319 74
rect -353 -74 -319 -58
rect -257 58 -223 74
rect -257 -74 -223 -58
rect -161 58 -127 74
rect -161 -74 -127 -58
rect -65 58 -31 74
rect -65 -74 -31 -58
rect 31 58 65 74
rect 31 -74 65 -58
rect 127 58 161 74
rect 127 -74 161 -58
rect 223 58 257 74
rect 223 -74 257 -58
rect 319 58 353 74
rect 319 -74 353 -58
rect 415 58 449 74
rect 415 -74 449 -58
rect 511 58 545 74
rect 511 -74 545 -58
rect 607 58 641 74
rect 607 -74 641 -58
rect 703 58 737 74
rect 703 -74 737 -58
rect -705 -151 -689 -117
rect -655 -151 -639 -117
rect 639 -151 655 -117
rect 689 -151 705 -117
rect -851 -219 -817 -157
rect 817 -219 851 -157
rect -851 -253 -755 -219
rect 755 -253 851 -219
<< viali >>
rect -593 117 -559 151
rect -497 117 -463 151
rect -401 117 -367 151
rect -305 117 -271 151
rect -209 117 -175 151
rect -113 117 -79 151
rect -17 117 17 151
rect 79 117 113 151
rect 175 117 209 151
rect 271 117 305 151
rect 367 117 401 151
rect 463 117 497 151
rect 559 117 593 151
rect -737 -58 -703 58
rect -641 -58 -607 58
rect -545 -58 -511 58
rect -449 -58 -415 58
rect -353 -58 -319 58
rect -257 -58 -223 58
rect -161 -58 -127 58
rect -65 -58 -31 58
rect 31 -58 65 58
rect 127 -58 161 58
rect 223 -58 257 58
rect 319 -58 353 58
rect 415 -58 449 58
rect 511 -58 545 58
rect 607 -58 641 58
rect 703 -58 737 58
rect -689 -151 -655 -117
rect 655 -151 689 -117
<< metal1 >>
rect -605 151 -547 157
rect -509 151 -451 157
rect -413 151 -355 157
rect -317 151 -259 157
rect -221 151 -163 157
rect -125 151 -67 157
rect -29 151 29 157
rect 67 151 125 157
rect 163 151 221 157
rect 259 151 317 157
rect 355 151 413 157
rect 451 151 509 157
rect 547 151 605 157
rect -609 117 -593 151
rect -559 117 -497 151
rect -463 117 -401 151
rect -367 117 -305 151
rect -271 117 -209 151
rect -175 117 -113 151
rect -79 117 -17 151
rect 17 117 79 151
rect 113 117 175 151
rect 209 117 271 151
rect 305 117 367 151
rect 401 117 463 151
rect 497 117 559 151
rect 593 117 609 151
rect -605 111 -547 117
rect -509 111 -451 117
rect -413 111 -355 117
rect -317 111 -259 117
rect -221 111 -163 117
rect -125 111 -67 117
rect -29 111 29 117
rect 67 111 125 117
rect 163 111 221 117
rect 259 111 317 117
rect 355 111 413 117
rect 451 111 509 117
rect 547 111 605 117
rect -752 66 -688 70
rect -752 14 -746 66
rect -694 14 -688 66
rect -752 6 -737 14
rect -743 -58 -737 6
rect -703 6 -688 14
rect -656 66 -592 70
rect -656 14 -650 66
rect -598 14 -592 66
rect -656 6 -641 14
rect -703 -58 -697 6
rect -743 -70 -697 -58
rect -647 -58 -641 6
rect -607 6 -592 14
rect -551 58 -505 70
rect -607 -58 -601 6
rect -551 -6 -545 58
rect -647 -70 -601 -58
rect -560 -12 -545 -6
rect -511 -6 -505 58
rect -464 66 -400 70
rect -464 14 -458 66
rect -406 14 -400 66
rect -464 6 -449 14
rect -511 -12 -496 -6
rect -560 -64 -554 -12
rect -502 -64 -496 -12
rect -560 -70 -496 -64
rect -455 -58 -449 6
rect -415 6 -400 14
rect -359 58 -313 70
rect -415 -58 -409 6
rect -359 -6 -353 58
rect -455 -70 -409 -58
rect -368 -12 -353 -6
rect -319 -6 -313 58
rect -272 66 -208 70
rect -272 14 -266 66
rect -214 14 -208 66
rect -272 6 -257 14
rect -319 -12 -304 -6
rect -368 -64 -362 -12
rect -310 -64 -304 -12
rect -368 -70 -304 -64
rect -263 -58 -257 6
rect -223 6 -208 14
rect -167 58 -121 70
rect -223 -58 -217 6
rect -167 -6 -161 58
rect -263 -70 -217 -58
rect -176 -12 -161 -6
rect -127 -6 -121 58
rect -80 66 -16 70
rect -80 14 -74 66
rect -22 14 -16 66
rect -80 6 -65 14
rect -127 -12 -112 -6
rect -176 -64 -170 -12
rect -118 -64 -112 -12
rect -176 -70 -112 -64
rect -71 -58 -65 6
rect -31 6 -16 14
rect 25 58 71 70
rect -31 -58 -25 6
rect 25 -6 31 58
rect -71 -70 -25 -58
rect 16 -12 31 -6
rect 65 -6 71 58
rect 112 66 176 70
rect 112 14 118 66
rect 170 14 176 66
rect 112 6 127 14
rect 65 -12 80 -6
rect 16 -64 22 -12
rect 74 -64 80 -12
rect 16 -70 80 -64
rect 121 -58 127 6
rect 161 6 176 14
rect 217 58 263 70
rect 161 -58 167 6
rect 217 -6 223 58
rect 121 -70 167 -58
rect 208 -12 223 -6
rect 257 -6 263 58
rect 304 66 368 70
rect 304 14 310 66
rect 362 14 368 66
rect 304 6 319 14
rect 257 -12 272 -6
rect 208 -64 214 -12
rect 266 -64 272 -12
rect 208 -70 272 -64
rect 313 -58 319 6
rect 353 6 368 14
rect 409 58 455 70
rect 353 -58 359 6
rect 409 -6 415 58
rect 313 -70 359 -58
rect 400 -12 415 -6
rect 449 -6 455 58
rect 496 66 560 70
rect 496 14 502 66
rect 554 14 560 66
rect 496 6 511 14
rect 449 -12 464 -6
rect 400 -64 406 -12
rect 458 -64 464 -12
rect 400 -70 464 -64
rect 505 -58 511 6
rect 545 6 560 14
rect 601 58 647 70
rect 545 -58 551 6
rect 601 -6 607 58
rect 505 -70 551 -58
rect 592 -12 607 -6
rect 641 -6 647 58
rect 688 66 752 70
rect 688 14 694 66
rect 746 14 752 66
rect 688 6 703 14
rect 641 -12 656 -6
rect 592 -64 598 -12
rect 650 -64 656 -12
rect 592 -70 656 -64
rect 697 -58 703 6
rect 737 6 752 14
rect 737 -58 743 6
rect 697 -70 743 -58
rect -701 -117 -643 -111
rect 643 -117 701 -111
rect -701 -151 -689 -117
rect -655 -151 655 -117
rect 689 -151 701 -117
rect -701 -157 -643 -151
rect 643 -157 701 -151
<< via1 >>
rect -746 58 -694 66
rect -746 14 -737 58
rect -737 14 -703 58
rect -703 14 -694 58
rect -650 58 -598 66
rect -650 14 -641 58
rect -641 14 -607 58
rect -607 14 -598 58
rect -458 58 -406 66
rect -458 14 -449 58
rect -449 14 -415 58
rect -415 14 -406 58
rect -554 -58 -545 -12
rect -545 -58 -511 -12
rect -511 -58 -502 -12
rect -554 -64 -502 -58
rect -266 58 -214 66
rect -266 14 -257 58
rect -257 14 -223 58
rect -223 14 -214 58
rect -362 -58 -353 -12
rect -353 -58 -319 -12
rect -319 -58 -310 -12
rect -362 -64 -310 -58
rect -74 58 -22 66
rect -74 14 -65 58
rect -65 14 -31 58
rect -31 14 -22 58
rect -170 -58 -161 -12
rect -161 -58 -127 -12
rect -127 -58 -118 -12
rect -170 -64 -118 -58
rect 118 58 170 66
rect 118 14 127 58
rect 127 14 161 58
rect 161 14 170 58
rect 22 -58 31 -12
rect 31 -58 65 -12
rect 65 -58 74 -12
rect 22 -64 74 -58
rect 310 58 362 66
rect 310 14 319 58
rect 319 14 353 58
rect 353 14 362 58
rect 214 -58 223 -12
rect 223 -58 257 -12
rect 257 -58 266 -12
rect 214 -64 266 -58
rect 502 58 554 66
rect 502 14 511 58
rect 511 14 545 58
rect 545 14 554 58
rect 406 -58 415 -12
rect 415 -58 449 -12
rect 449 -58 458 -12
rect 406 -64 458 -58
rect 694 58 746 66
rect 694 14 703 58
rect 703 14 737 58
rect 737 14 746 58
rect 598 -58 607 -12
rect 607 -58 641 -12
rect 641 -58 650 -12
rect 598 -64 650 -58
<< metal2 >>
rect -757 68 -587 77
rect -757 12 -748 68
rect -692 12 -652 68
rect -596 12 -587 68
rect -757 3 -587 12
rect -469 68 -395 77
rect -469 12 -460 68
rect -404 12 -395 68
rect -469 3 -395 12
rect -277 68 -203 77
rect -277 12 -268 68
rect -212 12 -203 68
rect -277 3 -203 12
rect -85 68 -11 77
rect -85 12 -76 68
rect -20 12 -11 68
rect -85 3 -11 12
rect 107 68 181 77
rect 107 12 116 68
rect 172 12 181 68
rect 107 3 181 12
rect 299 68 373 77
rect 299 12 308 68
rect 364 12 373 68
rect 299 3 373 12
rect 491 68 565 77
rect 491 12 500 68
rect 556 12 565 68
rect 491 3 565 12
rect 683 68 757 77
rect 683 12 692 68
rect 748 12 757 68
rect 683 3 757 12
rect -560 -12 -496 -6
rect -560 -64 -554 -12
rect -502 -36 -496 -12
rect -368 -12 -304 -6
rect -368 -36 -362 -12
rect -502 -64 -362 -36
rect -310 -36 -304 -12
rect -176 -12 -112 -6
rect -176 -36 -170 -12
rect -310 -64 -170 -36
rect -118 -36 -112 -12
rect 16 -12 80 -6
rect 16 -36 22 -12
rect -118 -64 22 -36
rect 74 -64 80 -12
rect -560 -70 80 -64
rect 208 -12 272 -6
rect 208 -64 214 -12
rect 266 -36 272 -12
rect 400 -12 464 -6
rect 400 -36 406 -12
rect 266 -64 406 -36
rect 458 -36 464 -12
rect 592 -12 656 -6
rect 592 -36 598 -12
rect 458 -64 598 -36
rect 650 -64 656 -12
rect 208 -70 656 -64
rect -257 -290 -223 -70
<< via2 >>
rect -748 66 -692 68
rect -748 14 -746 66
rect -746 14 -694 66
rect -694 14 -692 66
rect -748 12 -692 14
rect -652 66 -596 68
rect -652 14 -650 66
rect -650 14 -598 66
rect -598 14 -596 66
rect -652 12 -596 14
rect -460 66 -404 68
rect -460 14 -458 66
rect -458 14 -406 66
rect -406 14 -404 66
rect -460 12 -404 14
rect -268 66 -212 68
rect -268 14 -266 66
rect -266 14 -214 66
rect -214 14 -212 66
rect -268 12 -212 14
rect -76 66 -20 68
rect -76 14 -74 66
rect -74 14 -22 66
rect -22 14 -20 66
rect -76 12 -20 14
rect 116 66 172 68
rect 116 14 118 66
rect 118 14 170 66
rect 170 14 172 66
rect 116 12 172 14
rect 308 66 364 68
rect 308 14 310 66
rect 310 14 362 66
rect 362 14 364 66
rect 308 12 364 14
rect 500 66 556 68
rect 500 14 502 66
rect 502 14 554 66
rect 554 14 556 66
rect 500 12 556 14
rect 692 66 748 68
rect 692 14 694 66
rect 694 14 746 66
rect 746 14 748 66
rect 692 12 748 14
<< metal3 >>
rect -757 70 -587 77
rect -469 70 -395 77
rect -277 70 -203 77
rect -85 70 -11 77
rect 107 70 181 77
rect 299 70 373 77
rect 491 70 565 77
rect 683 70 757 77
rect -757 68 757 70
rect -757 12 -748 68
rect -692 12 -652 68
rect -596 12 -460 68
rect -404 12 -268 68
rect -212 12 -76 68
rect -20 12 116 68
rect 172 12 308 68
rect 364 12 500 68
rect 556 12 692 68
rect 748 12 757 68
rect -757 10 757 12
rect -757 3 -587 10
rect -469 3 -395 10
rect -277 3 -203 10
rect -85 3 -11 10
rect 107 3 181 10
rect 299 3 373 10
rect 491 3 565 10
rect 683 3 757 10
<< properties >>
string FIXED_BBOX -834 -236 834 236
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.7 l 0.15 m 1 nf 15 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
