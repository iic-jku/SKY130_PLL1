magic
tech sky130A
magscale 1 2
timestamp 1668153059
<< pwell >>
rect -455 -280 455 280
<< nmos >>
rect -255 -70 -225 70
rect -159 -70 -129 70
rect -63 -70 -33 70
rect 33 -70 63 70
rect 129 -70 159 70
rect 225 -70 255 70
<< ndiff >>
rect -317 58 -255 70
rect -317 -58 -305 58
rect -271 -58 -255 58
rect -317 -70 -255 -58
rect -225 58 -159 70
rect -225 -58 -209 58
rect -175 -58 -159 58
rect -225 -70 -159 -58
rect -129 58 -63 70
rect -129 -58 -113 58
rect -79 -58 -63 58
rect -129 -70 -63 -58
rect -33 58 33 70
rect -33 -58 -17 58
rect 17 -58 33 58
rect -33 -70 33 -58
rect 63 58 129 70
rect 63 -58 79 58
rect 113 -58 129 58
rect 63 -70 129 -58
rect 159 58 225 70
rect 159 -58 175 58
rect 209 -58 225 58
rect 159 -70 225 -58
rect 255 58 317 70
rect 255 -58 271 58
rect 305 0 317 58
rect 305 -58 318 0
rect 255 -70 318 -58
<< ndiffc >>
rect -305 -58 -271 58
rect -209 -58 -175 58
rect -113 -58 -79 58
rect -17 -58 17 58
rect 79 -58 113 58
rect 175 -58 209 58
rect 271 -58 305 58
<< psubdiff >>
rect -419 210 -323 244
rect 323 210 419 244
rect -419 148 -385 210
rect 385 148 419 210
rect -419 -210 -385 -148
rect 385 -210 419 -148
rect -419 -244 -323 -210
rect 323 -244 419 -210
<< psubdiffcont >>
rect -323 210 323 244
rect -419 -148 -385 148
rect 385 -148 419 148
rect -323 -244 323 -210
<< poly >>
rect -177 142 177 158
rect -177 108 -161 142
rect -127 108 -65 142
rect -31 108 31 142
rect 65 108 127 142
rect 161 108 177 142
rect -255 70 -225 96
rect -177 92 177 108
rect -159 70 -129 92
rect -63 70 -33 92
rect 33 70 63 92
rect 129 70 159 92
rect 225 70 255 96
rect -255 -92 -225 -70
rect -273 -108 -207 -92
rect -159 -96 -129 -70
rect -63 -96 -33 -70
rect 33 -96 63 -70
rect 129 -96 159 -70
rect 225 -92 255 -70
rect -273 -142 -257 -108
rect -223 -142 -207 -108
rect -273 -158 -207 -142
rect 207 -108 273 -92
rect 207 -142 223 -108
rect 257 -142 273 -108
rect 207 -158 273 -142
<< polycont >>
rect -161 108 -127 142
rect -65 108 -31 142
rect 31 108 65 142
rect 127 108 161 142
rect -257 -142 -223 -108
rect 223 -142 257 -108
<< locali >>
rect -419 210 -323 244
rect 323 210 419 244
rect -419 148 -385 210
rect 385 148 419 210
rect -177 108 -161 142
rect -127 108 -65 142
rect -31 108 31 142
rect 65 108 127 142
rect 161 108 177 142
rect -305 58 -271 74
rect -305 -74 -271 -58
rect -209 58 -175 74
rect -209 -74 -175 -58
rect -113 58 -79 74
rect -113 -74 -79 -58
rect -17 58 17 74
rect -17 -74 17 -58
rect 79 58 113 74
rect 79 -74 113 -58
rect 175 58 209 74
rect 175 -74 209 -58
rect 271 58 305 74
rect 271 -74 305 -58
rect -273 -142 -257 -108
rect -223 -142 -207 -108
rect 207 -142 223 -108
rect 257 -142 273 -108
rect -419 -210 -385 -148
rect 385 -210 419 -148
rect -419 -244 -323 -210
rect 323 -244 419 -210
<< viali >>
rect -161 108 -127 142
rect -65 108 -31 142
rect 31 108 65 142
rect 127 108 161 142
rect -305 -58 -271 58
rect -209 -58 -175 58
rect -113 -58 -79 58
rect -17 -58 17 58
rect 79 -58 113 58
rect 175 -58 209 58
rect 271 -58 305 58
rect -257 -142 -223 -108
rect 223 -142 257 -108
<< metal1 >>
rect -173 142 173 148
rect -173 108 -161 142
rect -127 108 -65 142
rect -31 108 31 142
rect 65 108 127 142
rect 161 108 173 142
rect -173 102 173 108
rect -311 58 -265 70
rect -311 0 -305 58
rect -317 -9 -305 0
rect -271 0 -265 58
rect -215 58 -169 70
rect -215 0 -209 58
rect -271 -9 -209 0
rect -175 0 -169 58
rect -125 61 -66 70
rect -125 9 -122 61
rect -70 28 -66 61
rect -23 58 23 70
rect -70 9 -67 28
rect -125 0 -113 9
rect -175 -9 -163 0
rect -317 -61 -314 -9
rect -262 -61 -218 -9
rect -166 -61 -163 -9
rect -317 -70 -163 -61
rect -119 -58 -113 0
rect -79 0 -67 9
rect -23 0 -17 58
rect -79 -58 -73 0
rect -119 -70 -73 -58
rect -29 -9 -17 0
rect 17 0 23 58
rect 67 61 125 70
rect 67 9 70 61
rect 122 9 125 61
rect 67 0 79 9
rect 17 -9 29 0
rect -29 -61 -26 -9
rect 26 -28 29 -9
rect 26 -61 30 -28
rect -29 -70 30 -61
rect 73 -58 79 0
rect 113 0 125 9
rect 169 58 215 70
rect 169 0 175 58
rect 113 -58 119 0
rect 73 -70 119 -58
rect 163 -9 175 0
rect 209 0 215 58
rect 265 58 311 70
rect 265 0 271 58
rect 209 -9 271 0
rect 305 0 311 58
rect 305 -9 318 0
rect 163 -61 166 -9
rect 218 -61 262 -9
rect 314 -61 318 -9
rect 163 -70 318 -61
rect -305 -102 -269 -70
rect 269 -102 305 -70
rect -305 -108 -211 -102
rect 211 -108 305 -102
rect -305 -142 -257 -108
rect -223 -142 -207 -108
rect 207 -142 223 -108
rect 257 -142 305 -108
rect -269 -148 -211 -142
rect 211 -148 269 -142
<< via1 >>
rect -122 58 -70 61
rect -122 9 -113 58
rect -113 9 -79 58
rect -79 9 -70 58
rect -314 -58 -305 -9
rect -305 -58 -271 -9
rect -271 -58 -262 -9
rect -314 -61 -262 -58
rect -218 -58 -209 -9
rect -209 -58 -175 -9
rect -175 -58 -166 -9
rect -218 -61 -166 -58
rect 70 58 122 61
rect 70 9 79 58
rect 79 9 113 58
rect 113 9 122 58
rect -26 -58 -17 -9
rect -17 -58 17 -9
rect 17 -58 26 -9
rect -26 -61 26 -58
rect 166 -58 175 -9
rect 175 -58 209 -9
rect 209 -58 218 -9
rect 166 -61 218 -58
rect 262 -58 271 -9
rect 271 -58 305 -9
rect 305 -58 314 -9
rect 262 -61 314 -58
<< metal2 >>
rect -125 61 125 70
rect -125 9 -122 61
rect -70 28 70 61
rect -70 9 -67 28
rect -125 0 -67 9
rect 67 9 70 28
rect 122 9 125 61
rect 67 0 125 9
rect -317 -9 -163 0
rect -317 -61 -314 -9
rect -262 -61 -218 -9
rect -166 -28 -163 -9
rect -29 -9 29 0
rect -29 -28 -26 -9
rect -166 -61 -26 -28
rect 26 -28 29 -9
rect 163 -9 318 0
rect 163 -28 166 -9
rect 26 -61 166 -28
rect 218 -61 262 -9
rect 314 -61 318 -9
rect -317 -70 318 -61
<< properties >>
string FIXED_BBOX -402 -227 402 227
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.7 l 0.150 m 1 nf 6 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
