magic
tech sky130A
magscale 1 2
timestamp 1660914963
<< locali >>
rect 2190 1934 2311 2104
rect 2140 1221 2203 1734
rect -970 -617 -800 -496
rect -600 -667 0 -604
rect 5068 -655 5668 -592
rect 5868 -605 6038 -484
rect 2781 -2998 2844 -2485
rect 2831 -3368 2952 -3198
<< metal1 >>
rect -1170 2104 6238 2304
rect -1170 -3368 -970 2104
rect -800 1734 5868 1934
rect -800 -2998 -600 1734
rect 2508 -135 2560 -129
rect 2508 -193 2560 -187
rect 2372 -416 2424 -410
rect 2372 -474 2424 -468
rect 2381 -790 2415 -474
rect 2372 -796 2424 -790
rect 2372 -854 2424 -848
rect 2517 -1071 2551 -193
rect 2644 -518 2696 -512
rect 2644 -576 2696 -570
rect 2653 -688 2687 -576
rect 2644 -694 2696 -688
rect 2644 -752 2696 -746
rect 2508 -1077 2560 -1071
rect 2508 -1135 2560 -1129
rect 5668 -2998 5868 1734
rect -800 -3198 5868 -2998
rect 6038 -3368 6238 2104
rect -1170 -3568 6238 -3368
<< via1 >>
rect 2508 -187 2560 -135
rect 2372 -468 2424 -416
rect 2372 -848 2424 -796
rect 2644 -570 2696 -518
rect 2644 -746 2696 -694
rect 2508 -1129 2560 -1077
<< metal2 >>
rect 1229 1295 1305 1305
rect 1229 1239 1239 1295
rect 1295 1239 1305 1295
rect 1229 1229 1305 1239
rect 2496 1293 2572 1303
rect 2496 1237 2506 1293
rect 2562 1282 2572 1293
rect 2562 1248 3818 1282
rect 2562 1237 2572 1248
rect 1250 1223 1284 1229
rect 2496 1227 2572 1237
rect 3784 1223 3818 1248
rect 1245 -37 1289 85
rect 2502 -187 2508 -135
rect 2560 -187 2566 -135
rect 2366 -468 2372 -416
rect 2424 -468 2430 -416
rect 2638 -570 2644 -518
rect 2696 -570 2702 -518
rect 1232 -604 1302 -597
rect 3766 -604 3836 -597
rect 1230 -660 1239 -604
rect 1295 -615 1304 -604
rect 3764 -615 3773 -604
rect 1295 -649 3773 -615
rect 1295 -660 1304 -649
rect 3764 -660 3773 -649
rect 3829 -660 3838 -604
rect 1232 -667 1302 -660
rect 3766 -667 3836 -660
rect 2638 -746 2644 -694
rect 2696 -746 2702 -694
rect 2366 -848 2372 -796
rect 2424 -848 2430 -796
rect 2502 -1086 2508 -1077
rect 2484 -1120 2508 -1086
rect 2502 -1129 2508 -1120
rect 2560 -1086 2566 -1077
rect 2560 -1120 2586 -1086
rect 2560 -1129 2566 -1120
rect 1250 -2512 1284 -2487
rect 2496 -2501 2572 -2491
rect 3784 -2493 3818 -2487
rect 2496 -2512 2506 -2501
rect 1250 -2546 2506 -2512
rect 2496 -2557 2506 -2546
rect 2562 -2557 2572 -2501
rect 2496 -2567 2572 -2557
rect 3763 -2503 3839 -2493
rect 3763 -2559 3773 -2503
rect 3829 -2559 3839 -2503
rect 3763 -2569 3839 -2559
<< via2 >>
rect 1239 1239 1295 1295
rect 2506 1237 2562 1293
rect 1239 -660 1295 -604
rect 3773 -660 3829 -604
rect 2506 -2557 2562 -2501
rect 3773 -2559 3829 -2503
<< metal3 >>
rect 1237 1311 1297 1342
rect 1223 1299 1311 1311
rect 1223 1235 1235 1299
rect 1299 1235 1311 1299
rect 1223 1223 1311 1235
rect 2490 1297 2578 1309
rect 2490 1233 2502 1297
rect 2566 1294 2578 1297
rect 2566 1234 2609 1294
rect 2566 1233 2578 1234
rect 2490 1221 2578 1233
rect -60 943 0 1003
rect 5068 943 5128 1003
rect -60 295 0 355
rect 5068 295 5128 355
rect 1223 73 1311 85
rect 1223 9 1235 73
rect 1299 9 1311 73
rect 1223 -3 1311 9
rect 2490 73 2578 85
rect 2490 9 2502 73
rect 2566 9 2578 73
rect 2490 -3 2578 9
rect 537 -140 597 -107
rect 528 -147 606 -140
rect 528 -211 535 -147
rect 599 -211 606 -147
rect 528 -218 606 -211
rect 528 -665 606 -658
rect 528 -729 535 -665
rect 599 -729 606 -665
rect 528 -736 606 -729
rect 537 -1157 597 -736
rect 834 -787 894 -107
rect 1237 -597 1297 -3
rect 1232 -604 1302 -597
rect 1232 -660 1239 -604
rect 1295 -660 1302 -604
rect 1639 -658 1699 -107
rect 1936 -269 1996 -107
rect 1927 -276 2005 -269
rect 1927 -340 1934 -276
rect 1998 -340 2005 -276
rect 1927 -347 2005 -340
rect 1232 -667 1302 -660
rect 1630 -665 1708 -658
rect 1630 -729 1637 -665
rect 1701 -729 1708 -665
rect 1630 -736 1708 -729
rect 825 -794 903 -787
rect 825 -858 832 -794
rect 896 -858 903 -794
rect 825 -865 903 -858
rect 1927 -794 2005 -787
rect 1927 -858 1934 -794
rect 1998 -858 2005 -794
rect 1927 -865 2005 -858
rect 1630 -924 1708 -917
rect 1630 -988 1637 -924
rect 1701 -988 1708 -924
rect 1630 -995 1708 -988
rect 825 -1053 903 -1046
rect 825 -1117 832 -1053
rect 896 -1117 903 -1053
rect 825 -1124 903 -1117
rect 834 -1157 894 -1124
rect 1639 -1157 1699 -995
rect 1936 -1157 1996 -865
rect 2504 -1261 2564 -3
rect 3072 -399 3132 -107
rect 3369 -140 3429 -107
rect 3360 -147 3438 -140
rect 3360 -211 3367 -147
rect 3431 -211 3438 -147
rect 3360 -218 3438 -211
rect 4174 -269 4234 -107
rect 4165 -276 4243 -269
rect 4165 -340 4172 -276
rect 4236 -340 4243 -276
rect 4165 -347 4243 -340
rect 3063 -406 3141 -399
rect 3063 -470 3070 -406
rect 3134 -470 3141 -406
rect 3063 -477 3141 -470
rect 3360 -406 3438 -399
rect 3360 -470 3367 -406
rect 3431 -470 3438 -406
rect 3360 -477 3438 -470
rect 3063 -1053 3141 -1046
rect 3063 -1117 3070 -1053
rect 3134 -1117 3141 -1053
rect 3063 -1124 3141 -1117
rect 3072 -1157 3132 -1124
rect 3369 -1157 3429 -477
rect 4471 -528 4531 -107
rect 4165 -535 4243 -528
rect 3766 -604 3836 -597
rect 3766 -660 3773 -604
rect 3829 -660 3836 -604
rect 4165 -599 4172 -535
rect 4236 -599 4243 -535
rect 4165 -606 4243 -599
rect 4462 -535 4540 -528
rect 4462 -599 4469 -535
rect 4533 -599 4540 -535
rect 4462 -606 4540 -599
rect 3766 -667 3836 -660
rect 3771 -1261 3831 -667
rect 4174 -1157 4234 -606
rect 4462 -924 4540 -917
rect 4462 -988 4469 -924
rect 4533 -988 4540 -924
rect 4462 -995 4540 -988
rect 4471 -1157 4531 -995
rect 2490 -1273 2578 -1261
rect 2490 -1337 2502 -1273
rect 2566 -1337 2578 -1273
rect 2490 -1349 2578 -1337
rect 3757 -1273 3845 -1261
rect 3757 -1337 3769 -1273
rect 3833 -1337 3845 -1273
rect 3757 -1349 3845 -1337
rect -60 -1619 0 -1559
rect 5068 -1619 5128 -1559
rect -60 -2267 0 -2207
rect 5068 -2267 5128 -2207
rect 2490 -2497 2578 -2485
rect 2490 -2498 2502 -2497
rect 2459 -2558 2502 -2498
rect 2490 -2561 2502 -2558
rect 2566 -2561 2578 -2497
rect 2490 -2573 2578 -2561
rect 3757 -2499 3845 -2487
rect 3757 -2563 3769 -2499
rect 3833 -2563 3845 -2499
rect 3757 -2575 3845 -2563
rect 3771 -2606 3831 -2575
<< via3 >>
rect 1235 1295 1299 1299
rect 1235 1239 1239 1295
rect 1239 1239 1295 1295
rect 1295 1239 1299 1295
rect 1235 1235 1299 1239
rect 2502 1293 2566 1297
rect 2502 1237 2506 1293
rect 2506 1237 2562 1293
rect 2562 1237 2566 1293
rect 2502 1233 2566 1237
rect 1235 9 1299 73
rect 2502 9 2566 73
rect 535 -211 599 -147
rect 535 -729 599 -665
rect 1934 -340 1998 -276
rect 1637 -729 1701 -665
rect 832 -858 896 -794
rect 1934 -858 1998 -794
rect 1637 -988 1701 -924
rect 832 -1117 896 -1053
rect 3367 -211 3431 -147
rect 4172 -340 4236 -276
rect 3070 -470 3134 -406
rect 3367 -470 3431 -406
rect 3070 -1117 3134 -1053
rect 4172 -599 4236 -535
rect 4469 -599 4533 -535
rect 4469 -988 4533 -924
rect 2502 -1337 2566 -1273
rect 3769 -1337 3833 -1273
rect 2502 -2501 2566 -2497
rect 2502 -2557 2506 -2501
rect 2506 -2557 2562 -2501
rect 2562 -2557 2566 -2501
rect 2502 -2561 2566 -2557
rect 3769 -2503 3833 -2499
rect 3769 -2559 3773 -2503
rect 3773 -2559 3829 -2503
rect 3829 -2559 3833 -2503
rect 3769 -2563 3833 -2559
<< metal4 >>
rect 1223 1299 1311 1311
rect 686 1221 746 1281
rect 1223 1235 1235 1299
rect 1299 1235 1311 1299
rect 2490 1297 2578 1309
rect 1223 1223 1311 1235
rect 1237 85 1297 1223
rect 1788 1221 1848 1281
rect 2490 1233 2502 1297
rect 2566 1233 2578 1297
rect 2490 1221 2578 1233
rect 3220 1221 3280 1281
rect 4322 1221 4382 1281
rect 2504 85 2564 1221
rect 1223 73 1311 85
rect 1223 9 1235 73
rect 1299 9 1311 73
rect 1223 -3 1311 9
rect 2490 73 2578 85
rect 2490 9 2502 73
rect 2566 9 2578 73
rect 2490 -3 2578 9
rect 528 -147 606 -140
rect 528 -149 535 -147
rect 0 -209 535 -149
rect 528 -211 535 -209
rect 599 -149 606 -147
rect 3360 -147 3438 -140
rect 3360 -149 3367 -147
rect 599 -209 3367 -149
rect 599 -211 606 -209
rect 528 -218 606 -211
rect 3360 -211 3367 -209
rect 3431 -149 3438 -147
rect 3431 -209 5068 -149
rect 3431 -211 3438 -209
rect 3360 -218 3438 -211
rect 1927 -276 2005 -269
rect 1927 -278 1934 -276
rect 0 -338 1934 -278
rect 1927 -340 1934 -338
rect 1998 -278 2005 -276
rect 4165 -276 4243 -269
rect 4165 -278 4172 -276
rect 1998 -338 4172 -278
rect 1998 -340 2005 -338
rect 1927 -347 2005 -340
rect 4165 -340 4172 -338
rect 4236 -278 4243 -276
rect 4236 -338 5068 -278
rect 4236 -340 4243 -338
rect 4165 -347 4243 -340
rect 3063 -406 3141 -399
rect 3063 -408 3070 -406
rect 0 -468 3070 -408
rect 3063 -470 3070 -468
rect 3134 -408 3141 -406
rect 3360 -406 3438 -399
rect 3360 -408 3367 -406
rect 3134 -468 3367 -408
rect 3134 -470 3141 -468
rect 3063 -477 3141 -470
rect 3360 -470 3367 -468
rect 3431 -408 3438 -406
rect 3431 -468 5068 -408
rect 3431 -470 3438 -468
rect 3360 -477 3438 -470
rect 4165 -535 4243 -528
rect 4165 -537 4172 -535
rect 0 -597 4172 -537
rect 4165 -599 4172 -597
rect 4236 -537 4243 -535
rect 4462 -535 4540 -528
rect 4462 -537 4469 -535
rect 4236 -597 4469 -537
rect 4236 -599 4243 -597
rect 4165 -606 4243 -599
rect 4462 -599 4469 -597
rect 4533 -537 4540 -535
rect 4533 -597 5068 -537
rect 4533 -599 4540 -597
rect 4462 -606 4540 -599
rect 528 -665 606 -658
rect 528 -667 535 -665
rect 0 -727 535 -667
rect 528 -729 535 -727
rect 599 -667 606 -665
rect 1630 -665 1708 -658
rect 1630 -667 1637 -665
rect 599 -727 1637 -667
rect 599 -729 606 -727
rect 528 -736 606 -729
rect 1630 -729 1637 -727
rect 1701 -667 1708 -665
rect 1701 -727 5068 -667
rect 1701 -729 1708 -727
rect 1630 -736 1708 -729
rect 825 -794 903 -787
rect 825 -796 832 -794
rect 0 -856 832 -796
rect 825 -858 832 -856
rect 896 -796 903 -794
rect 1927 -794 2005 -787
rect 1927 -796 1934 -794
rect 896 -856 1934 -796
rect 896 -858 903 -856
rect 825 -865 903 -858
rect 1927 -858 1934 -856
rect 1998 -796 2005 -794
rect 1998 -856 5068 -796
rect 1998 -858 2005 -856
rect 1927 -865 2005 -858
rect 1630 -924 1708 -917
rect 1630 -926 1637 -924
rect 0 -986 1637 -926
rect 1630 -988 1637 -986
rect 1701 -926 1708 -924
rect 4462 -924 4540 -917
rect 4462 -926 4469 -924
rect 1701 -986 4469 -926
rect 1701 -988 1708 -986
rect 1630 -995 1708 -988
rect 4462 -988 4469 -986
rect 4533 -926 4540 -924
rect 4533 -986 5068 -926
rect 4533 -988 4540 -986
rect 4462 -995 4540 -988
rect 825 -1053 903 -1046
rect 825 -1055 832 -1053
rect 0 -1115 832 -1055
rect 825 -1117 832 -1115
rect 896 -1055 903 -1053
rect 3063 -1053 3141 -1046
rect 3063 -1055 3070 -1053
rect 896 -1115 3070 -1055
rect 896 -1117 903 -1115
rect 825 -1124 903 -1117
rect 3063 -1117 3070 -1115
rect 3134 -1055 3141 -1053
rect 3134 -1115 5068 -1055
rect 3134 -1117 3141 -1115
rect 3063 -1124 3141 -1117
rect 2490 -1273 2578 -1261
rect 2490 -1337 2502 -1273
rect 2566 -1337 2578 -1273
rect 2490 -1349 2578 -1337
rect 3757 -1273 3845 -1261
rect 3757 -1337 3769 -1273
rect 3833 -1337 3845 -1273
rect 3757 -1349 3845 -1337
rect 2504 -2485 2564 -1349
rect 686 -2545 746 -2485
rect 1788 -2545 1848 -2485
rect 2490 -2497 2578 -2485
rect 2490 -2561 2502 -2497
rect 2566 -2561 2578 -2497
rect 3220 -2545 3280 -2485
rect 3771 -2487 3831 -1349
rect 3757 -2499 3845 -2487
rect 2490 -2573 2578 -2561
rect 3757 -2563 3769 -2499
rect 3833 -2563 3845 -2499
rect 4322 -2545 4382 -2485
rect 3757 -2575 3845 -2563
use delay_cell_4  delay_cell_4_0
timestamp 1660732324
transform 1 0 865 0 1 138
box -865 -735 1669 1085
use delay_cell_4  delay_cell_4_1
timestamp 1660732324
transform -1 0 4203 0 1 138
box -865 -735 1669 1085
use delay_cell_4  delay_cell_4_2
timestamp 1660732324
transform -1 0 4203 0 -1 -1402
box -865 -735 1669 1085
use delay_cell_4  delay_cell_4_3
timestamp 1660732324
transform 1 0 865 0 -1 -1402
box -865 -735 1669 1085
<< labels >>
rlabel metal3 5068 943 5128 1003 0 vdd
rlabel metal3 5068 -2267 5128 -2207 0 vdd
rlabel metal3 5068 -1619 5128 -1559 0 vss
rlabel metal3 5068 295 5128 355 0 vss
rlabel metal2 3784 1223 3818 1282 0 vb1
rlabel metal4 1223 1223 1311 1311 0 vb2
rlabel metal4 528 -218 606 -140 0 out1
rlabel metal4 1927 -347 2005 -269 0 out2
rlabel metal4 3063 -477 3141 -399 7 out3
rlabel metal4 4462 -606 4540 -528 0 out4
rlabel metal4 4462 -995 4540 -917 0 out5
rlabel metal4 3063 -1124 3141 -1046 3 out6
rlabel metal4 1927 -865 2005 -787 5 out7
rlabel metal4 528 -736 606 -658 0 out8
rlabel metal1 2653 -649 2687 -615 7 b0
rlabel metal1 2517 -649 2551 -615 0 b1
rlabel metal1 2381 -649 2415 -615 0 b2
rlabel metal4 686 1221 746 1281 0 inv1
rlabel metal4 1788 1221 1848 1281 0 inv2
rlabel metal4 3220 1221 3280 1281 0 inv3
rlabel metal4 4322 1221 4382 1281 6 inv4
rlabel metal4 4322 -2545 4382 -2485 7 inv5
rlabel metal4 3220 -2545 3280 -2485 3 inv6
rlabel metal4 1788 -2545 1848 -2485 4 inv7
rlabel metal4 686 -2545 746 -2485 7 inv8
<< end >>
