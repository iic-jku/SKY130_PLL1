magic
tech sky130A
magscale 1 2
timestamp 1668153059
<< pwell >>
rect -8631 -2369 8631 2369
<< psubdiff >>
rect -8595 2299 -8499 2333
rect 8499 2299 8595 2333
rect -8595 2237 -8561 2299
rect 8561 2237 8595 2299
rect -8595 -2299 -8561 -2237
rect 8561 -2299 8595 -2237
rect -8595 -2333 -8499 -2299
rect 8499 -2333 8595 -2299
<< psubdiffcont >>
rect -8499 2299 8499 2333
rect -8595 -2237 -8561 2237
rect 8561 -2237 8595 2237
rect -8499 -2333 8499 -2299
<< xpolycontact >>
rect -8465 1771 -7895 2203
rect -8465 -2203 -7895 -1771
rect -7647 1771 -7077 2203
rect -7647 -2203 -7077 -1771
rect -6829 1771 -6259 2203
rect -6829 -2203 -6259 -1771
rect -6011 1771 -5441 2203
rect -6011 -2203 -5441 -1771
rect -5193 1771 -4623 2203
rect -5193 -2203 -4623 -1771
rect -4375 1771 -3805 2203
rect -4375 -2203 -3805 -1771
rect -3557 1771 -2987 2203
rect -3557 -2203 -2987 -1771
rect -2739 1771 -2169 2203
rect -2739 -2203 -2169 -1771
rect -1921 1771 -1351 2203
rect -1921 -2203 -1351 -1771
rect -1103 1771 -533 2203
rect -1103 -2203 -533 -1771
rect -285 1771 285 2203
rect -285 -2203 285 -1771
rect 533 1771 1103 2203
rect 533 -2203 1103 -1771
rect 1351 1771 1921 2203
rect 1351 -2203 1921 -1771
rect 2169 1771 2739 2203
rect 2169 -2203 2739 -1771
rect 2987 1771 3557 2203
rect 2987 -2203 3557 -1771
rect 3805 1771 4375 2203
rect 3805 -2203 4375 -1771
rect 4623 1771 5193 2203
rect 4623 -2203 5193 -1771
rect 5441 1771 6011 2203
rect 5441 -2203 6011 -1771
rect 6259 1771 6829 2203
rect 6259 -2203 6829 -1771
rect 7077 1771 7647 2203
rect 7077 -2203 7647 -1771
rect 7895 1771 8465 2203
rect 7895 -2203 8465 -1771
<< ppolyres >>
rect -8465 -1771 -7895 1771
rect -7647 -1771 -7077 1771
rect -6829 -1771 -6259 1771
rect -6011 -1771 -5441 1771
rect -5193 -1771 -4623 1771
rect -4375 -1771 -3805 1771
rect -3557 -1771 -2987 1771
rect -2739 -1771 -2169 1771
rect -1921 -1771 -1351 1771
rect -1103 -1771 -533 1771
rect -285 -1771 285 1771
rect 533 -1771 1103 1771
rect 1351 -1771 1921 1771
rect 2169 -1771 2739 1771
rect 2987 -1771 3557 1771
rect 3805 -1771 4375 1771
rect 4623 -1771 5193 1771
rect 5441 -1771 6011 1771
rect 6259 -1771 6829 1771
rect 7077 -1771 7647 1771
rect 7895 -1771 8465 1771
<< locali >>
rect -8595 2299 -8499 2333
rect 8499 2299 8595 2333
rect -8595 2237 -8561 2299
rect 8561 2237 8595 2299
rect -8595 -2299 -8561 -2237
rect 8561 -2299 8595 -2237
rect -8595 -2333 -8499 -2299
rect 8499 -2333 8595 -2299
<< viali >>
rect -8449 1788 -7911 2185
rect -7631 1788 -7093 2185
rect -6813 1788 -6275 2185
rect -5995 1788 -5457 2185
rect -5177 1788 -4639 2185
rect -4359 1788 -3821 2185
rect -3541 1788 -3003 2185
rect -2723 1788 -2185 2185
rect -1905 1788 -1367 2185
rect -1087 1788 -549 2185
rect -269 1788 269 2185
rect 549 1788 1087 2185
rect 1367 1788 1905 2185
rect 2185 1788 2723 2185
rect 3003 1788 3541 2185
rect 3821 1788 4359 2185
rect 4639 1788 5177 2185
rect 5457 1788 5995 2185
rect 6275 1788 6813 2185
rect 7093 1788 7631 2185
rect 7911 1788 8449 2185
rect -8449 -2185 -7911 -1788
rect -7631 -2185 -7093 -1788
rect -6813 -2185 -6275 -1788
rect -5995 -2185 -5457 -1788
rect -5177 -2185 -4639 -1788
rect -4359 -2185 -3821 -1788
rect -3541 -2185 -3003 -1788
rect -2723 -2185 -2185 -1788
rect -1905 -2185 -1367 -1788
rect -1087 -2185 -549 -1788
rect -269 -2185 269 -1788
rect 549 -2185 1087 -1788
rect 1367 -2185 1905 -1788
rect 2185 -2185 2723 -1788
rect 3003 -2185 3541 -1788
rect 3821 -2185 4359 -1788
rect 4639 -2185 5177 -1788
rect 5457 -2185 5995 -1788
rect 6275 -2185 6813 -1788
rect 7093 -2185 7631 -1788
rect 7911 -2185 8449 -1788
<< metal1 >>
rect -8461 2185 -7899 2191
rect -8461 1788 -8449 2185
rect -7911 1788 -7899 2185
rect -8461 1782 -7899 1788
rect -7643 2185 -7081 2191
rect -7643 1788 -7631 2185
rect -7093 1788 -7081 2185
rect -7643 1782 -7081 1788
rect -6825 2185 -6263 2191
rect -6825 1788 -6813 2185
rect -6275 1788 -6263 2185
rect -6825 1782 -6263 1788
rect -6007 2185 -5445 2191
rect -6007 1788 -5995 2185
rect -5457 1788 -5445 2185
rect -6007 1782 -5445 1788
rect -5189 2185 -4627 2191
rect -5189 1788 -5177 2185
rect -4639 1788 -4627 2185
rect -5189 1782 -4627 1788
rect -4371 2185 -3809 2191
rect -4371 1788 -4359 2185
rect -3821 1788 -3809 2185
rect -4371 1782 -3809 1788
rect -3553 2185 -2991 2191
rect -3553 1788 -3541 2185
rect -3003 1788 -2991 2185
rect -3553 1782 -2991 1788
rect -2735 2185 -2173 2191
rect -2735 1788 -2723 2185
rect -2185 1788 -2173 2185
rect -2735 1782 -2173 1788
rect -1917 2185 -1355 2191
rect -1917 1788 -1905 2185
rect -1367 1788 -1355 2185
rect -1917 1782 -1355 1788
rect -1099 2185 -537 2191
rect -1099 1788 -1087 2185
rect -549 1788 -537 2185
rect -1099 1782 -537 1788
rect -281 2185 281 2191
rect -281 1788 -269 2185
rect 269 1788 281 2185
rect -281 1782 281 1788
rect 537 2185 1099 2191
rect 537 1788 549 2185
rect 1087 1788 1099 2185
rect 537 1782 1099 1788
rect 1355 2185 1917 2191
rect 1355 1788 1367 2185
rect 1905 1788 1917 2185
rect 1355 1782 1917 1788
rect 2173 2185 2735 2191
rect 2173 1788 2185 2185
rect 2723 1788 2735 2185
rect 2173 1782 2735 1788
rect 2991 2185 3553 2191
rect 2991 1788 3003 2185
rect 3541 1788 3553 2185
rect 2991 1782 3553 1788
rect 3809 2185 4371 2191
rect 3809 1788 3821 2185
rect 4359 1788 4371 2185
rect 3809 1782 4371 1788
rect 4627 2185 5189 2191
rect 4627 1788 4639 2185
rect 5177 1788 5189 2185
rect 4627 1782 5189 1788
rect 5445 2185 6007 2191
rect 5445 1788 5457 2185
rect 5995 1788 6007 2185
rect 5445 1782 6007 1788
rect 6263 2185 6825 2191
rect 6263 1788 6275 2185
rect 6813 1788 6825 2185
rect 6263 1782 6825 1788
rect 7081 2185 7643 2191
rect 7081 1788 7093 2185
rect 7631 1788 7643 2185
rect 7081 1782 7643 1788
rect 7899 2185 8461 2191
rect 7899 1788 7911 2185
rect 8449 1788 8461 2185
rect 7899 1782 8461 1788
rect -8461 -1788 -7899 -1782
rect -8461 -2185 -8449 -1788
rect -7911 -2185 -7899 -1788
rect -8461 -2191 -7899 -2185
rect -7643 -1788 -7081 -1782
rect -7643 -2185 -7631 -1788
rect -7093 -2185 -7081 -1788
rect -7643 -2191 -7081 -2185
rect -6825 -1788 -6263 -1782
rect -6825 -2185 -6813 -1788
rect -6275 -2185 -6263 -1788
rect -6825 -2191 -6263 -2185
rect -6007 -1788 -5445 -1782
rect -6007 -2185 -5995 -1788
rect -5457 -2185 -5445 -1788
rect -6007 -2191 -5445 -2185
rect -5189 -1788 -4627 -1782
rect -5189 -2185 -5177 -1788
rect -4639 -2185 -4627 -1788
rect -5189 -2191 -4627 -2185
rect -4371 -1788 -3809 -1782
rect -4371 -2185 -4359 -1788
rect -3821 -2185 -3809 -1788
rect -4371 -2191 -3809 -2185
rect -3553 -1788 -2991 -1782
rect -3553 -2185 -3541 -1788
rect -3003 -2185 -2991 -1788
rect -3553 -2191 -2991 -2185
rect -2735 -1788 -2173 -1782
rect -2735 -2185 -2723 -1788
rect -2185 -2185 -2173 -1788
rect -2735 -2191 -2173 -2185
rect -1917 -1788 -1355 -1782
rect -1917 -2185 -1905 -1788
rect -1367 -2185 -1355 -1788
rect -1917 -2191 -1355 -2185
rect -1099 -1788 -537 -1782
rect -1099 -2185 -1087 -1788
rect -549 -2185 -537 -1788
rect -1099 -2191 -537 -2185
rect -281 -1788 281 -1782
rect -281 -2185 -269 -1788
rect 269 -2185 281 -1788
rect -281 -2191 281 -2185
rect 537 -1788 1099 -1782
rect 537 -2185 549 -1788
rect 1087 -2185 1099 -1788
rect 537 -2191 1099 -2185
rect 1355 -1788 1917 -1782
rect 1355 -2185 1367 -1788
rect 1905 -2185 1917 -1788
rect 1355 -2191 1917 -2185
rect 2173 -1788 2735 -1782
rect 2173 -2185 2185 -1788
rect 2723 -2185 2735 -1788
rect 2173 -2191 2735 -2185
rect 2991 -1788 3553 -1782
rect 2991 -2185 3003 -1788
rect 3541 -2185 3553 -1788
rect 2991 -2191 3553 -2185
rect 3809 -1788 4371 -1782
rect 3809 -2185 3821 -1788
rect 4359 -2185 4371 -1788
rect 3809 -2191 4371 -2185
rect 4627 -1788 5189 -1782
rect 4627 -2185 4639 -1788
rect 5177 -2185 5189 -1788
rect 4627 -2191 5189 -2185
rect 5445 -1788 6007 -1782
rect 5445 -2185 5457 -1788
rect 5995 -2185 6007 -1788
rect 5445 -2191 6007 -2185
rect 6263 -1788 6825 -1782
rect 6263 -2185 6275 -1788
rect 6813 -2185 6825 -1788
rect 6263 -2191 6825 -2185
rect 7081 -1788 7643 -1782
rect 7081 -2185 7093 -1788
rect 7631 -2185 7643 -1788
rect 7081 -2191 7643 -2185
rect 7899 -1788 8461 -1782
rect 7899 -2185 7911 -1788
rect 8449 -2185 8461 -1788
rect 7899 -2191 8461 -2185
<< res2p85 >>
rect -8467 -1773 -7893 1773
rect -7649 -1773 -7075 1773
rect -6831 -1773 -6257 1773
rect -6013 -1773 -5439 1773
rect -5195 -1773 -4621 1773
rect -4377 -1773 -3803 1773
rect -3559 -1773 -2985 1773
rect -2741 -1773 -2167 1773
rect -1923 -1773 -1349 1773
rect -1105 -1773 -531 1773
rect -287 -1773 287 1773
rect 531 -1773 1105 1773
rect 1349 -1773 1923 1773
rect 2167 -1773 2741 1773
rect 2985 -1773 3559 1773
rect 3803 -1773 4377 1773
rect 4621 -1773 5195 1773
rect 5439 -1773 6013 1773
rect 6257 -1773 6831 1773
rect 7075 -1773 7649 1773
rect 7893 -1773 8467 1773
<< properties >>
string FIXED_BBOX -8578 -2316 8578 2316
string gencell sky130_fd_pr__res_high_po_2p85
string library sky130
string parameters w 2.850 l 17.71 m 1 nx 21 wmin 2.850 lmin 0.50 rho 319.8 val 2.0k dummy 0 dw 0.0 term 19.188 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} full_metal 1 wmax 2.850 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
